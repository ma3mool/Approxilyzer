
module decode_unit ( instruction, o_rd, o_rd_type, o_rd_valid, o_rd2, 
        o_rd2_type, o_rd2_valid, o_rs1, o_rs1_type, o_rs1_valid, o_rs2, 
        o_rs2_type, o_rs2_valid, o_rs3, o_rs3_type, o_rs3_valid, o_rs4, 
        o_rs4_type, o_rs4_valid, o_m_type, o_m_futype, o_m_opcode, 
        o_m_branch_type, o_m_imm, o_m_ccshift, o_m_access_size, o_m_flags, 
        o_fail );
  input [31:0] instruction;
  output [5:0] o_rd;
  output [3:0] o_rd_type;
  output [5:0] o_rd2;
  output [3:0] o_rd2_type;
  output [5:0] o_rs1;
  output [3:0] o_rs1_type;
  output [5:0] o_rs2;
  output [3:0] o_rs2_type;
  output [5:0] o_rs3;
  output [3:0] o_rs3_type;
  output [5:0] o_rs4;
  output [3:0] o_rs4_type;
  output [2:0] o_m_type;
  output [3:0] o_m_futype;
  output [8:0] o_m_opcode;
  output [3:0] o_m_branch_type;
  output [63:0] o_m_imm;
  output [7:0] o_m_ccshift;
  output [7:0] o_m_access_size;
  output [7:0] o_m_flags;
  output o_rd_valid, o_rd2_valid, o_rs1_valid, o_rs2_valid, o_rs3_valid,
         o_rs4_valid, o_fail;
  wire   n_Logic0_, o_rs2_4_, o_rs2_3_, o_rs2_2_, o_rs2_1_, o_rs4_valid, N5185,
         N5186, N5187, N5188, N5189, n250, n360, n378, n379, n387, n388, n390,
         n395, n399, n400, n409, n410, n412, n415, n416, n424, n425, n441,
         n457, n470, n472, n475, n488, n528, n535, n587, n590, n591, n593,
         n594, n595, n599, n631, n633, n644, n647, n671, n674, n679, n681,
         n834, n835, n840, n874, n885, n919, n922, n930, n990, n992, n1084,
         n1093, n1094, n1095, n1128, n1133, n1137, n1139, n1161, n1229, n1230,
         n1231, n1375, n1383, n1395, n1405, n1407, n1422, n1442, n1443, n1544,
         n1549, n1550, n673, r944_carry_2_, r944_carry_3_, r944_carry_4_,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, o_m_imm_38_, o_m_imm_40_, o_m_imm_42_, o_m_imm_44_,
         o_m_imm_48_, o_m_imm_52_, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, o_m_access_size_6_, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989;
  assign o_m_flags[0] = n_Logic0_;
  assign o_m_flags[7] = n_Logic0_;
  assign o_m_access_size[5] = n_Logic0_;
  assign o_m_ccshift[0] = n_Logic0_;
  assign o_m_ccshift[3] = n_Logic0_;
  assign o_m_ccshift[4] = n_Logic0_;
  assign o_m_ccshift[5] = n_Logic0_;
  assign o_m_ccshift[6] = n_Logic0_;
  assign o_m_ccshift[7] = n_Logic0_;
  assign o_rs4_type[0] = n_Logic0_;
  assign o_rs4_type[1] = n_Logic0_;
  assign o_rs4_type[3] = n_Logic0_;
  assign o_rs2_type[3] = n_Logic0_;
  assign o_rs1_type[3] = n_Logic0_;
  assign o_rs2[4] = o_rs2_4_;
  assign o_rs2_4_ = instruction[4];
  assign o_rs2[3] = o_rs2_3_;
  assign o_rs2_3_ = instruction[3];
  assign o_rs2[2] = o_rs2_2_;
  assign o_rs2_2_ = instruction[2];
  assign o_rs2[1] = o_rs2_1_;
  assign o_rs2_1_ = instruction[1];
  assign o_rs4_type[2] = o_rs4_valid;
  assign o_m_imm[56] = o_m_imm_38_;
  assign o_m_imm[51] = o_m_imm_38_;
  assign o_m_imm[43] = o_m_imm_38_;
  assign o_m_imm[36] = o_m_imm_38_;
  assign o_m_imm[38] = o_m_imm_38_;
  assign o_m_imm[35] = o_m_imm_40_;
  assign o_m_imm[53] = o_m_imm_40_;
  assign o_m_imm[45] = o_m_imm_40_;
  assign o_m_imm[34] = o_m_imm_40_;
  assign o_m_imm[40] = o_m_imm_40_;
  assign o_m_imm[59] = o_m_imm_42_;
  assign o_m_imm[50] = o_m_imm_42_;
  assign o_m_imm[55] = o_m_imm_42_;
  assign o_m_imm[60] = o_m_imm_42_;
  assign o_m_imm[32] = o_m_imm_42_;
  assign o_m_imm[42] = o_m_imm_42_;
  assign o_m_imm[63] = o_m_imm_44_;
  assign o_m_imm[57] = o_m_imm_44_;
  assign o_m_imm[58] = o_m_imm_44_;
  assign o_m_imm[33] = o_m_imm_44_;
  assign o_m_imm[44] = o_m_imm_44_;
  assign o_m_imm[46] = o_m_imm_48_;
  assign o_m_imm[39] = o_m_imm_48_;
  assign o_m_imm[61] = o_m_imm_48_;
  assign o_m_imm[54] = o_m_imm_48_;
  assign o_m_imm[37] = o_m_imm_48_;
  assign o_m_imm[48] = o_m_imm_48_;
  assign o_m_imm[62] = o_m_imm_52_;
  assign o_m_imm[47] = o_m_imm_52_;
  assign o_m_imm[49] = o_m_imm_52_;
  assign o_m_imm[41] = o_m_imm_52_;
  assign o_m_imm[52] = o_m_imm_52_;
  assign o_rs3_type[3] = o_m_access_size_6_;
  assign o_m_access_size[6] = o_m_access_size_6_;

  HDNOR2D1 U705 ( .A1(instruction[13]), .A2(instruction[12]), .Z(n1422) );
  HDNAN2D1 U242 ( .A1(instruction[8]), .A2(n2972), .Z(n441) );
  HDNOR3D1 U378 ( .A1(n2981), .A2(n2980), .A3(instruction[8]), .Z(n591) );
  HDNAN3D1 U373 ( .A1(instruction[5]), .A2(instruction[8]), .A3(n2980), .Z(
        n647) );
  HDNAN2D1 U370 ( .A1(n647), .A2(n992), .Z(n874) );
  HDNOR2D1 U369 ( .A1(n1407), .A2(n874), .Z(n1405) );
  HDNOR2D1 U813 ( .A1(o_rs2_1_), .A2(instruction[0]), .Z(n1443) );
  HDNOR2D1 U88 ( .A1(n2975), .A2(n2974), .Z(n681) );
  HDNAN2D1 U746 ( .A1(instruction[7]), .A2(n1230), .Z(n930) );
  HDNAN2D1 U273 ( .A1(n2984), .A2(n2979), .Z(n1139) );
  HDNAN2D1 U272 ( .A1(n2985), .A2(n1139), .Z(n1231) );
  HDNOR3D1 U246 ( .A1(instruction[5]), .A2(n2979), .A3(n2980), .Z(n990) );
  HDNOR2D1 U255 ( .A1(n2971), .A2(n2975), .Z(n644) );
  HDNOR2D1 U50 ( .A1(n528), .A2(n1732), .Z(o_rs1[5]) );
  HDNOR2D1 U149 ( .A1(n2976), .A2(n834), .Z(n593) );
  HDNAN2D1 U81 ( .A1(n647), .A2(n2989), .Z(n590) );
  HDAOI211D1 U1337 ( .A1(n2968), .A2(n2967), .B(n488), .C(n919), .Z(n1375) );
  HDOAI21D1 U1330 ( .A1(n1375), .A2(n1732), .B(n475), .Z(o_m_futype[3]) );
  HDOAI211D1 U1474 ( .A1(n2980), .A2(n2979), .B(n2989), .C(n595), .Z(n1549) );
  HDNOR4D1 U1164 ( .A1(n2966), .A2(n2964), .A3(n472), .A4(n1095), .Z(n1093) );
  HDNAN2D1 U184 ( .A1(instruction[7]), .A2(n2979), .Z(n1084) );
  HDOR2D1 U1381 ( .A1(o_rd2_type[3]), .A2(o_rd2_type[2]), .Z(o_m_flags[4]) );
  HDAOI211D1 U974 ( .A1(n2968), .A2(n415), .B(n593), .C(n594), .Z(n587) );
  HDAOI31D1 U906 ( .A1(n399), .A2(n400), .A3(n2961), .B(n1732), .Z(
        o_rs2_type[2]) );
  HDOAI211D1 U900 ( .A1(instruction[11]), .A2(n360), .B(n378), .C(n379), .Z(
        o_rs3[0]) );
  HDNOR2D2 U828 ( .A1(instruction[11]), .A2(instruction[10]), .Z(n1544) );
  HDNAN2DL U374 ( .A1(n2983), .A2(n2985), .Z(n1407) );
  HDAOI211D1 U989 ( .A1(n2968), .A2(n2973), .B(n2964), .C(n593), .Z(n631) );
  HDNOR2D2 U381 ( .A1(n2960), .A2(n2959), .Z(n671) );
  HDOAI22D1 U1187 ( .A1(n2965), .A2(n2987), .B1(n1137), .B2(n835), .Z(n1128)
         );
  HDOAI211DL U1468 ( .A1(n2988), .A2(n1383), .B(n2977), .C(n470), .Z(n1550) );
  HDAOI31D1 U1165 ( .A1(n457), .A2(n992), .A3(n679), .B(n2987), .Z(n1095) );
  HDNAN2D1 U72 ( .A1(n633), .A2(n2985), .Z(n395) );
  HDOAI211D1 U924 ( .A1(n2971), .A2(n409), .B(instruction[12]), .C(n2969), .Z(
        n412) );
  HDAOI21D1 U910 ( .A1(n416), .A2(n415), .B(n2966), .Z(n410) );
  HDAOI21D1 U934 ( .A1(n2963), .A2(n2962), .B(n1732), .Z(o_rs1_type[2]) );
  HDADHALFD1 r944_U1_1_2 ( .A(instruction[27]), .B(r944_carry_2_), .CO(
        r944_carry_3_), .S(N5186) );
  HDADHALFD1 r944_U1_1_4 ( .A(instruction[29]), .B(r944_carry_4_), .CO(N5189), 
        .S(N5188) );
  HDADHALFD1 r944_U1_1_3 ( .A(instruction[28]), .B(r944_carry_3_), .CO(
        r944_carry_4_), .S(N5187) );
  HDADHALFD1 r944_U1_1_1 ( .A(instruction[26]), .B(instruction[25]), .CO(
        r944_carry_2_), .S(N5185) );
  HDNAN4D1 U1483 ( .A1(n1801), .A2(n2502), .A3(n2676), .A4(n2733), .Z(n1910)
         );
  HDNOR2D1 U1484 ( .A1(n1686), .A2(n2732), .Z(n1800) );
  HDNAN2D1 U1485 ( .A1(n2001), .A2(n2162), .Z(n2029) );
  HDNAN2D1 U1486 ( .A1(n2932), .A2(n2931), .Z(n2936) );
  HDAND2D1 U1487 ( .A1(n1927), .A2(n1928), .Z(n1942) );
  HDINVBD2 U1488 ( .A(n2018), .Z(n1831) );
  HDINVBD2 U1489 ( .A(n2777), .Z(n2658) );
  HDNOR2D1 U1490 ( .A1(n2524), .A2(n1715), .Z(n2478) );
  HDINVD8 U1491 ( .A(instruction[21]), .Z(n2374) );
  HDINVD2 U1492 ( .A(n2934), .Z(n2941) );
  HDINVD2 U1493 ( .A(instruction[13]), .Z(n2977) );
  HDAND2D1 U1494 ( .A1(n2760), .A2(n1599), .Z(n2849) );
  HDINVD12 U1495 ( .A(instruction[27]), .Z(n2948) );
  HDINVD1 U1496 ( .A(n1731), .Z(n1869) );
  HDNOR2D1 U1497 ( .A1(n2560), .A2(instruction[14]), .Z(n1842) );
  HDAND2D1 U1498 ( .A1(n1823), .A2(n2323), .Z(n2505) );
  HDAND2D1 U1499 ( .A1(n2969), .A2(instruction[12]), .Z(n2158) );
  HDINVD1 U1500 ( .A(n2508), .Z(n1821) );
  HDNOR2D1 U1501 ( .A1(n1951), .A2(instruction[24]), .Z(n1822) );
  HDNOR2D1 U1502 ( .A1(n1889), .A2(n2934), .Z(n1913) );
  HDNAN3D1 U1503 ( .A1(n1887), .A2(instruction[13]), .A3(n2738), .Z(n1891) );
  HDNOR3D1 U1504 ( .A1(n1910), .A2(n1912), .A3(n1617), .Z(n1914) );
  HDINVD1 U1505 ( .A(n1913), .Z(n1729) );
  HDINVD1 U1506 ( .A(n1868), .Z(n2256) );
  HDNOR2D6 U1507 ( .A1(n1774), .A2(instruction[19]), .Z(n2189) );
  HDNAN2D1 U1508 ( .A1(n2906), .A2(n2063), .Z(n2851) );
  HDINVD1 U1509 ( .A(n1873), .Z(n1704) );
  HDNAN3D1 U1510 ( .A1(n2399), .A2(n1947), .A3(n1161), .Z(n1796) );
  HDINVD1 U1511 ( .A(n1395), .Z(n2176) );
  HDNAN2D2 U1512 ( .A1(n2323), .A2(n2018), .Z(n2655) );
  HDINVD1 U1513 ( .A(n2860), .Z(n2632) );
  HDNAN2D1 U1514 ( .A1(n2322), .A2(n1865), .Z(n2418) );
  HDINVD2 U1515 ( .A(n2650), .Z(n2676) );
  HDNOR2D1 U1516 ( .A1(n2901), .A2(n2100), .Z(n2802) );
  HDNAN2D2 U1517 ( .A1(n1731), .A2(n2018), .Z(n2659) );
  HDAND2D1 U1518 ( .A1(n2973), .A2(instruction[7]), .Z(n2713) );
  HDNAN2D2 U1519 ( .A1(n1888), .A2(n2018), .Z(n2450) );
  HDINVBD2 U1520 ( .A(n2004), .Z(n2548) );
  HDNAN4D1 U1521 ( .A1(n2214), .A2(n2658), .A3(n2952), .A4(n2029), .Z(n2002)
         );
  HDNOR2D1 U1522 ( .A1(n2309), .A2(instruction[25]), .Z(n2760) );
  HDINVD1 U1523 ( .A(instruction[30]), .Z(n1892) );
  HDINVD1 U1524 ( .A(n2500), .Z(n1812) );
  HDINVD1 U1525 ( .A(n1657), .Z(n1604) );
  HDINVD1 U1526 ( .A(n2936), .Z(n1605) );
  HDINVD1 U1527 ( .A(n2865), .Z(n2916) );
  HDNOR4D1 U1528 ( .A1(n1781), .A2(n1780), .A3(n1919), .A4(n1779), .Z(n1829)
         );
  HDNOR2D1 U1529 ( .A1(n1732), .A2(n2399), .Z(n1927) );
  HDNOR2D1 U1530 ( .A1(n1922), .A2(n1736), .Z(n1908) );
  HDINVD2 U1531 ( .A(n1936), .Z(n1926) );
  HDNOR2D2 U1532 ( .A1(n2533), .A2(n2497), .Z(n1936) );
  HDINVBD2 U1533 ( .A(instruction[10]), .Z(n2978) );
  HDINVD2 U1534 ( .A(instruction[11]), .Z(n2064) );
  HDAND2D1 U1535 ( .A1(n1967), .A2(n1602), .Z(n1965) );
  HDAND4D1 U1536 ( .A1(n1974), .A2(n1723), .A3(n1973), .A4(n1972), .Z(n1615)
         );
  HDNOR2D1 U1537 ( .A1(n2578), .A2(n2934), .Z(n2770) );
  HDNOR2D1 U1538 ( .A1(n2486), .A2(n2038), .Z(n1832) );
  HDINVD2 U1539 ( .A(n1688), .Z(n2492) );
  HDNOR2D1 U1540 ( .A1(n1796), .A2(n2176), .Z(n2968) );
  HDINVD1 U1541 ( .A(n2655), .Z(n2499) );
  HDINVD2 U1542 ( .A(n2603), .Z(n2567) );
  HDNOR2D1 U1543 ( .A1(n1835), .A2(n1688), .Z(n2586) );
  HDINVD1 U1544 ( .A(n2633), .Z(n1852) );
  HDNAN3D1 U1545 ( .A1(n1686), .A2(n2501), .A3(n1888), .Z(n2601) );
  HDINVD1 U1546 ( .A(n2859), .Z(n2628) );
  HDNAN2D1 U1547 ( .A1(n2305), .A2(n2601), .Z(n2634) );
  HDINVD1 U1548 ( .A(n2533), .Z(n2637) );
  HDOA31DL U1549 ( .A1(n2976), .A2(n2799), .A3(n2319), .B(n2800), .Z(n2664) );
  HDINVD2 U1550 ( .A(n2323), .Z(n2679) );
  HDINVD1 U1551 ( .A(n2687), .Z(n2693) );
  HDINVD1 U1552 ( .A(n388), .Z(n2799) );
  HDINVBD2 U1553 ( .A(n2987), .Z(n2723) );
  HDAOI21M20DL U1554 ( .A1(n2922), .A2(n2925), .B(n2930), .Z(n2743) );
  HDINVD1 U1555 ( .A(instruction[0]), .Z(n2746) );
  HDINVD1 U1556 ( .A(instruction[15]), .Z(n2809) );
  HDINVD4 U1557 ( .A(instruction[17]), .Z(n2811) );
  HDINVD2 U1558 ( .A(instruction[18]), .Z(n2812) );
  HDNOR3D1 U1559 ( .A1(n2372), .A2(n2040), .A3(n2834), .Z(n2816) );
  HDINVD1 U1560 ( .A(n1732), .Z(n1735) );
  HDNAN2D1 U1561 ( .A1(n1607), .A2(n1609), .Z(n1656) );
  HDNAN3D1 U1562 ( .A1(n1604), .A2(n1605), .A3(n1606), .Z(n1607) );
  HDINVD1 U1563 ( .A(n2933), .Z(n1606) );
  HDINVD8 U1564 ( .A(instruction[28]), .Z(n2951) );
  HDINVD1 U1565 ( .A(n2497), .Z(n1600) );
  HDAOI211D1 U1566 ( .A1(n2942), .A2(n1609), .B(n2941), .C(n1599), .Z(n2953)
         );
  HDOAI21M20DL U1567 ( .A1(n2449), .A2(n2448), .B(n1609), .Z(n2457) );
  HDAO22DL U1568 ( .A1(n2849), .A2(N5189), .B1(n2848), .B2(n1735), .Z(o_rd2[5]) );
  HDOA211DL U1569 ( .A1(n2394), .A2(n2798), .B(n2422), .C(n2398), .Z(n1558) );
  HDAND3D1 U1570 ( .A1(n2411), .A2(n1616), .A3(n1558), .Z(n2307) );
  HDNAN2M1D1 U1571 ( .A1(n2113), .A2(n595), .Z(n409) );
  HDNOR2M1D1 U1572 ( .A1(n2331), .A2(n2666), .Z(n1559) );
  HDNAN4D1 U1573 ( .A1(n2511), .A2(n2477), .A3(n2459), .A4(n1559), .Z(n2371)
         );
  HDAOI211D1 U1574 ( .A1(n2446), .A2(n2447), .B(n2441), .C(n2445), .Z(n1560)
         );
  HDOA211DL U1575 ( .A1(n2444), .A2(n2443), .B(n2442), .C(n1560), .Z(n2448) );
  HDAOI32D1 U1576 ( .A1(n671), .A2(n2491), .A3(n2468), .B1(n2852), .B2(n2491), 
        .Z(n1561) );
  HDNOR3D1 U1577 ( .A1(n2470), .A2(n2469), .A3(n1561), .Z(n2473) );
  HDOAI21D1 U1578 ( .A1(n395), .A2(n599), .B(n2355), .Z(n400) );
  HDAOI21M20D1 U1579 ( .A1(instruction[25]), .A2(n1990), .B(n2213), .Z(n1995)
         );
  HDNAN3M1D1 U1580 ( .A1(n488), .A2(n2450), .A3(n2271), .Z(n2272) );
  HDNAN3D1 U1581 ( .A1(n2482), .A2(n2464), .A3(n2463), .Z(n1562) );
  HDNOR4D1 U1582 ( .A1(n2650), .A2(n2834), .A3(n2760), .A4(n1562), .Z(n2477)
         );
  HDNOR3M1D4 U1583 ( .A1(n1731), .A2(n1685), .A3(n2934), .Z(n2876) );
  HDNOR4M1D1 U1584 ( .A1(n2382), .A2(n2329), .A3(n2666), .A4(n1627), .Z(n1563)
         );
  HDNAN4D1 U1585 ( .A1(n2330), .A2(n2422), .A3(n2583), .A4(n1563), .Z(n1626)
         );
  HDNAN2M1D1 U1586 ( .A1(n2597), .A2(n2506), .Z(n2471) );
  HDOAI21D1 U1587 ( .A1(instruction[13]), .A2(n1829), .B(n2520), .Z(n1564) );
  HDNAN2D1 U1588 ( .A1(n1564), .A2(n1599), .Z(n390) );
  HDAO211DL U1589 ( .A1(n674), .A2(n2723), .B(n2721), .C(n2722), .Z(n1565) );
  HDINVDL U1590 ( .A(n2724), .Z(n1566) );
  HDOAI211D1 U1591 ( .A1(n2725), .A2(n2988), .B(n470), .C(n1566), .Z(n1567) );
  HDNOR4D1 U1592 ( .A1(n472), .A2(n2726), .A3(n1565), .A4(n1567), .Z(n2729) );
  HDNOR2M1D1 U1593 ( .A1(n2836), .A2(o_m_flags[3]), .Z(n2843) );
  HDOAI22D1 U1594 ( .A1(n1947), .A2(n2098), .B1(n2086), .B2(n2113), .Z(n1568)
         );
  HDNOR3M1D1 U1595 ( .A1(n1422), .A2(n2969), .A3(n1568), .Z(n2742) );
  HDNAN2M1D1 U1596 ( .A1(n2042), .A2(n2346), .Z(n2021) );
  HDNAN3D1 U1597 ( .A1(n2309), .A2(n2464), .A3(n2764), .Z(n1569) );
  HDOAI31D1 U1598 ( .A1(n2478), .A2(n2087), .A3(n1569), .B(instruction[10]), 
        .Z(n1921) );
  HDNOR3M1D1 U1599 ( .A1(n2550), .A2(n2030), .A3(n2146), .Z(n2032) );
  HDNAN4M1D1 U1600 ( .A1(n2371), .A2(n2476), .A3(n2376), .A4(n2451), .Z(n2381)
         );
  HDNAN2D1 U1601 ( .A1(n2655), .A2(n2493), .Z(n1570) );
  HDNOR4D1 U1602 ( .A1(n2494), .A2(n2648), .A3(n2920), .A4(n1570), .Z(n2677)
         );
  HDAOI21M20D1 U1603 ( .A1(n1836), .A2(n1867), .B(n1736), .Z(o_m_flags[2]) );
  HDAOI22D1 U1604 ( .A1(n2355), .A2(n2799), .B1(n2977), .B2(n1830), .Z(n1571)
         );
  HDAND4D1 U1605 ( .A1(n2530), .A2(n2882), .A3(n2961), .A4(n1571), .Z(n1572)
         );
  HDOAI21D1 U1606 ( .A1(n1732), .A2(n1572), .B(n390), .Z(o_rs2_valid) );
  HDINVDL U1607 ( .A(instruction[9]), .Z(n1573) );
  HDAO33DL U1608 ( .A1(n1573), .A2(instruction[5]), .A3(n1161), .B1(
        instruction[9]), .B2(n1544), .B3(n2176), .Z(n1809) );
  HDNAN2M1D1 U1609 ( .A1(n2213), .A2(n1601), .Z(n2148) );
  HDNAN3M1D1 U1610 ( .A1(n2373), .A2(n2511), .A3(n2251), .Z(n2329) );
  HDNAN2M1D1 U1611 ( .A1(n1845), .A2(n2310), .Z(n2626) );
  HDNOR2M1D1 U1612 ( .A1(n1770), .A2(n1687), .Z(n2372) );
  HDNAN3D1 U1613 ( .A1(n2598), .A2(n2596), .A3(n2597), .Z(n1574) );
  HDOAI31M10D1 U1614 ( .A1(n2615), .A2(n2599), .A3(n1574), .B(n2859), .Z(n2600) );
  HDNAN4DL U1615 ( .A1(n2763), .A2(n2764), .A3(n2818), .A4(n2765), .Z(n1575)
         );
  HDAOI31D1 U1616 ( .A1(n2767), .A2(n2769), .A3(n2768), .B(n1732), .Z(n1576)
         );
  HDAOI211D1 U1617 ( .A1(n1599), .A2(n1575), .B(n2770), .C(n1576), .Z(n2782)
         );
  HDAOI21M20DL U1618 ( .A1(n1829), .A2(n2977), .B(n1833), .Z(n1577) );
  HDNAN3D1 U1619 ( .A1(instruction[13]), .A2(n1830), .A3(n1734), .Z(n1578) );
  HDOAI211D1 U1620 ( .A1(n1737), .A2(n1577), .B(n2868), .C(n1578), .Z(
        o_m_flags[1]) );
  HDNAN2D1 U1621 ( .A1(n1863), .A2(n1719), .Z(n1579) );
  HDOAI211D1 U1622 ( .A1(n2583), .A2(n1866), .B(n2738), .C(n1579), .Z(n1580)
         );
  HDNOR3D1 U1623 ( .A1(n2041), .A2(n2252), .A3(n1580), .Z(n1581) );
  HDAOI31D1 U1624 ( .A1(n2264), .A2(n2130), .A3(n1581), .B(n1736), .Z(
        o_m_access_size[3]) );
  HDAOI211D1 U1625 ( .A1(n2723), .A2(n395), .B(n2711), .C(n2710), .Z(n1582) );
  HDAOI21M20DL U1626 ( .A1(n2929), .A2(n1582), .B(n2758), .Z(n1583) );
  HDOAI22M10D1 U1627 ( .A1(n2717), .A2(n2716), .B1(n1732), .B2(n1583), .Z(
        o_rs2_type[0]) );
  HDOAI211D1 U1628 ( .A1(instruction[8]), .A2(n2755), .B(n1644), .C(n2468), 
        .Z(n1584) );
  HDNOR2M1D1 U1629 ( .A1(n388), .A2(n1584), .Z(n1645) );
  HDNAN2M1D1 U1630 ( .A1(n2966), .A2(n2396), .Z(n2314) );
  HDNOR2M1D1 U1631 ( .A1(n2245), .A2(n2213), .Z(n2222) );
  HDNAN4M1D1 U1632 ( .A1(o_rs2_2_), .A2(n1443), .A3(n2977), .A4(n2716), .Z(
        n2423) );
  HDNOR2M1D1 U1633 ( .A1(n2560), .A2(n2561), .Z(n2627) );
  HDNOR3M1D1 U1634 ( .A1(n2759), .A2(n2761), .A3(n2760), .Z(n2765) );
  HDNOR3M1D1 U1635 ( .A1(n2727), .A2(n2085), .A3(n595), .Z(n2773) );
  HDAOI31D1 U1636 ( .A1(n2767), .A2(n1898), .A3(n2918), .B(n1732), .Z(n1585)
         );
  HDNOR2D1 U1637 ( .A1(n1915), .A2(n1585), .Z(n1897) );
  HDAND2D1 U1638 ( .A1(n1967), .A2(n1964), .Z(n1955) );
  HDOAI21M10D1 U1639 ( .A1(n2443), .A2(n2664), .B(n1609), .Z(n360) );
  HDNOR2M1D1 U1640 ( .A1(n2959), .A2(n2927), .Z(n2711) );
  HDNAN3M1D1 U1641 ( .A1(n2737), .A2(n2931), .A3(n2738), .Z(n2808) );
  HDNAN3D1 U1642 ( .A1(n2435), .A2(n2673), .A3(n2582), .Z(n1586) );
  HDNAN4D1 U1643 ( .A1(n1864), .A2(n2817), .A3(n2023), .A4(n2044), .Z(n1587)
         );
  HDAOI211D1 U1644 ( .A1(n2258), .A2(n2139), .B(n1586), .C(n1587), .Z(n1588)
         );
  HDNOR2D1 U1645 ( .A1(n1588), .A2(n1737), .Z(o_m_access_size[2]) );
  HDNOR3D1 U1646 ( .A1(n2870), .A2(n2020), .A3(n2087), .Z(n1589) );
  HDAOI21D1 U1647 ( .A1(n2641), .A2(n1589), .B(n1736), .Z(o_m_access_size[7])
         );
  HDOA211DL U1648 ( .A1(n425), .A2(n424), .B(instruction[0]), .C(n1735), .Z(
        o_rs2[5]) );
  HDNAN2M1D1 U1649 ( .A1(n2861), .A2(n1854), .Z(n1590) );
  HDOAI21M20DL U1650 ( .A1(n1590), .A2(n1609), .B(n2832), .Z(o_rd2_type[2]) );
  HDINVBD4 U1651 ( .A(n2231), .Z(n2944) );
  HDINVBD2 U1652 ( .A(n1599), .Z(n1736) );
  HDINVBD4 U1653 ( .A(n250), .Z(n1599) );
  HDNAN2D1 U1654 ( .A1(n1974), .A2(n1673), .Z(n1591) );
  HDNOR2D2 U1655 ( .A1(n2749), .A2(n2864), .Z(n1592) );
  HDNOR2D2 U1656 ( .A1(n2862), .A2(n1593), .Z(n1876) );
  HDINVD1 U1657 ( .A(n1592), .Z(n1593) );
  HDINVD4 U1658 ( .A(n2327), .Z(n1873) );
  HDINVD4 U1659 ( .A(n1966), .Z(n1967) );
  HDAND3D2 U1660 ( .A1(n2482), .A2(n2464), .A3(n2463), .Z(n1596) );
  HDNAN2D1 U1661 ( .A1(instruction[31]), .A2(instruction[30]), .Z(n250) );
  HDOR2D1 U1662 ( .A1(n2928), .A2(n673), .Z(n1594) );
  HDINVD1 U1663 ( .A(n1719), .Z(n1720) );
  HDAND2D1 U1664 ( .A1(n2732), .A2(n2376), .Z(n1595) );
  HDAND3D1 U1665 ( .A1(n2529), .A2(n2530), .A3(n2571), .Z(n1597) );
  HDINVD4 U1666 ( .A(instruction[12]), .Z(n2399) );
  HDOR2D1 U1667 ( .A1(n1768), .A2(n1769), .Z(n1598) );
  HDNAN2D1 U1668 ( .A1(n1653), .A2(n1600), .Z(o_rd[0]) );
  HDNOR4D2 U1669 ( .A1(n2808), .A2(n1732), .A3(n2807), .A4(n2806), .Z(n2813)
         );
  HDOAI211DL U1670 ( .A1(n2339), .A2(n1704), .B(n1628), .C(n1629), .Z(n1625)
         );
  HDINVD1 U1671 ( .A(n2849), .Z(n2828) );
  HDNAN2D1 U1672 ( .A1(n1953), .A2(n1952), .Z(n1971) );
  HDNAN2M1D1 U1673 ( .A1(n2770), .A2(n1937), .Z(n2533) );
  HDINVD1 U1674 ( .A(n1732), .Z(n1733) );
  HDOAI21D1 U1675 ( .A1(instruction[31]), .A2(n2377), .B(n1600), .Z(n1954) );
  HDINVD1 U1676 ( .A(n1968), .Z(n1969) );
  HDNOR2D4 U1677 ( .A1(n1892), .A2(instruction[31]), .Z(n2497) );
  HDNOR2D6 U1678 ( .A1(n1752), .A2(instruction[23]), .Z(n2323) );
  HDINVD1 U1679 ( .A(n1908), .Z(n1918) );
  HDOAI211DL U1680 ( .A1(n2825), .A2(n1732), .B(n2824), .C(n2828), .Z(
        o_rd2_valid) );
  HDOAI211DL U1681 ( .A1(n2690), .A2(n2934), .B(n2689), .C(n2688), .Z(o_rs3[2]) );
  HDINVD4 U1682 ( .A(n2876), .Z(n2868) );
  HDNAN2D1 U1683 ( .A1(n2967), .A2(n416), .Z(n2397) );
  HDOA22M20D1 U1684 ( .A1(n2176), .A2(n2787), .B1(n1645), .B2(n2927), .Z(n1641) );
  HDAND3D1 U1685 ( .A1(n2627), .A2(n2626), .A3(n2625), .Z(n2629) );
  HDINVBD2 U1686 ( .A(n1725), .Z(n2777) );
  HDOAI22D1 U1687 ( .A1(n2034), .A2(n2679), .B1(n2234), .B2(n1704), .Z(n2035)
         );
  HDINVD1 U1688 ( .A(n1970), .Z(n1602) );
  HDAOI21D1 U1689 ( .A1(n2679), .A2(n2377), .B(n2934), .Z(n2646) );
  HDINVD2 U1690 ( .A(n1599), .Z(n1737) );
  HDINVD12 U1691 ( .A(n1609), .Z(n1732) );
  HDNAN2DL U1692 ( .A1(n2678), .A2(instruction[21]), .Z(n2680) );
  HDINVD4 U1693 ( .A(instruction[29]), .Z(n2952) );
  HDNOR3D2 U1694 ( .A1(n2943), .A2(instruction[28]), .A3(instruction[27]), .Z(
        n2030) );
  HDBUFD1 U1695 ( .A(n2030), .Z(n1697) );
  HDAND2D4 U1696 ( .A1(n1777), .A2(n1951), .Z(n2257) );
  HDNAN2DL U1697 ( .A1(n2001), .A2(n2161), .Z(n1601) );
  HDNOR2D2 U1698 ( .A1(n2979), .A2(n885), .Z(n1133) );
  HDNAN2D1 U1699 ( .A1(n2704), .A2(n390), .Z(n2717) );
  HDINVD4 U1700 ( .A(n2893), .Z(n1700) );
  HDINVD4 U1701 ( .A(n2509), .Z(n1714) );
  HDOA21M20D1 U1702 ( .A1(n2301), .A2(n1609), .B(n1600), .Z(n2302) );
  HDNOR2D2 U1703 ( .A1(n1807), .A2(instruction[9]), .Z(n1759) );
  HDNAN3D2 U1704 ( .A1(n1760), .A2(n1759), .A3(n2113), .Z(n399) );
  HDINVD2 U1705 ( .A(n1897), .Z(n1893) );
  HDNAN2M1D1 U1706 ( .A1(n2509), .A2(n2696), .Z(n1725) );
  HDINVBD4 U1707 ( .A(n1715), .Z(n2265) );
  HDNAN2M1D2 U1708 ( .A1(n1620), .A2(n2719), .Z(n2721) );
  HDBUFD8 U1709 ( .A(n2777), .Z(n1686) );
  HDOA21D1 U1710 ( .A1(n2912), .A2(n2911), .B(n2955), .Z(n1603) );
  HDNAN2D1 U1711 ( .A1(n1603), .A2(n2910), .Z(o_rd_type[1]) );
  HDAND2D2 U1712 ( .A1(instruction[27]), .A2(instruction[28]), .Z(n2210) );
  HDNAN3D2 U1713 ( .A1(n1991), .A2(n2244), .A3(n2245), .Z(n1994) );
  HDOAI21M20D1 U1714 ( .A1(n2972), .A2(n2883), .B(n2882), .Z(n2884) );
  HDNOR3D2 U1715 ( .A1(n2504), .A2(n2864), .A3(n2503), .Z(n2919) );
  HDNOR2D1 U1716 ( .A1(n1591), .A2(n1970), .Z(n1716) );
  HDNAN2D1 U1717 ( .A1(n1597), .A2(n2531), .Z(n2532) );
  HDNOR2D6 U1718 ( .A1(n2810), .A2(instruction[15]), .Z(n2543) );
  HDBUFBD4 U1719 ( .A(n2338), .Z(n1688) );
  HDNAN2D6 U1720 ( .A1(n2210), .A2(n2162), .Z(n2245) );
  HDINVD2 U1721 ( .A(n1999), .Z(n2009) );
  HDNOR2D1 U1722 ( .A1(n2171), .A2(n2632), .Z(n2645) );
  HDINVD2 U1723 ( .A(n1759), .Z(n2086) );
  HDNOR3D2 U1724 ( .A1(n1659), .A2(n1660), .A3(n1594), .Z(n1658) );
  HDINVD2 U1725 ( .A(n2607), .Z(n2320) );
  HDNOR3D4 U1726 ( .A1(n2085), .A2(n1806), .A3(n1741), .Z(n2607) );
  HDNAN2D2 U1727 ( .A1(n1876), .A2(n1595), .Z(n1928) );
  HDNOR2D2 U1728 ( .A1(n2871), .A2(n1598), .Z(n2731) );
  HDAOI21M20D1 U1729 ( .A1(n1928), .A2(n2506), .B(n1732), .Z(n1920) );
  HDNAN2M1D2 U1730 ( .A1(n2964), .A2(n1661), .Z(n1659) );
  HDNAN3D1 U1731 ( .A1(n2158), .A2(n387), .A3(n1644), .Z(n1642) );
  HDOA21M20D2 U1732 ( .A1(n1890), .A2(n2977), .B(n1672), .Z(n1922) );
  HDNOR2D2 U1733 ( .A1(n2679), .A2(n1868), .Z(n2859) );
  HDNAN2D4 U1734 ( .A1(n2492), .A2(n1823), .Z(n2435) );
  HDAND2D2 U1735 ( .A1(n2827), .A2(n1879), .Z(n2458) );
  HDOAI211D1 U1736 ( .A1(n1701), .A2(n2912), .B(n1600), .C(n2891), .Z(
        o_rd_type[0]) );
  HDINVD32 U1737 ( .A(instruction[5]), .Z(n2982) );
  HDNOR2D6 U1738 ( .A1(n2982), .A2(instruction[6]), .Z(n2973) );
  HDNAN2D4 U1739 ( .A1(n2713), .A2(n2979), .Z(n2985) );
  HDAO21D2 U1740 ( .A1(n1922), .A2(n1921), .B(n250), .Z(n1673) );
  HDAND2D2 U1741 ( .A1(n2336), .A2(n2696), .Z(n2339) );
  HDINVD8 U1742 ( .A(instruction[25]), .Z(n2696) );
  HDNAN4D1 U1743 ( .A1(n2919), .A2(n2918), .A3(n2917), .A4(n1665), .Z(n1662)
         );
  HDINVD8 U1744 ( .A(n1700), .Z(n1701) );
  HDNAN4D1 U1745 ( .A1(n2307), .A2(n2269), .A3(n2268), .A4(n2267), .Z(n2273)
         );
  HDNOR2D6 U1746 ( .A1(n2579), .A2(n2243), .Z(n2789) );
  HDOAI21M20D2 U1747 ( .A1(n1839), .A2(instruction[18]), .B(n2055), .Z(n2119)
         );
  HDINVD8 U1748 ( .A(n1714), .Z(n1715) );
  HDAND3DL U1749 ( .A1(n1698), .A2(n1825), .A3(n1824), .Z(n1722) );
  HDNAN2DL U1750 ( .A1(n2257), .A2(n2018), .Z(n2121) );
  HDNOR2D6 U1751 ( .A1(n1743), .A2(instruction[20]), .Z(n2018) );
  HDNOR2DL U1752 ( .A1(n2980), .A2(n387), .Z(n673) );
  HDINVD2 U1753 ( .A(n2210), .Z(n1986) );
  HDOAI211DL U1754 ( .A1(n1756), .A2(n1715), .B(n2874), .C(n1755), .Z(n1757)
         );
  HDINVDL U1755 ( .A(n2624), .Z(n1717) );
  HDAOI22DL U1756 ( .A1(n1863), .A2(n1715), .B1(n2192), .B2(instruction[25]), 
        .Z(n1825) );
  HDOR2D2 U1757 ( .A1(n1715), .A2(n2696), .Z(n2617) );
  HDNAN4D2 U1758 ( .A1(n1761), .A2(n1701), .A3(n2399), .A4(n2948), .Z(n2935)
         );
  HDNAN2D2 U1759 ( .A1(instruction[25]), .A2(instruction[26]), .Z(n2949) );
  HDBUFD8 U1760 ( .A(n2949), .Z(n1689) );
  HDINVD4 U1761 ( .A(n2881), .Z(n2929) );
  HDNOR2D4 U1762 ( .A1(n1861), .A2(n2243), .Z(n2739) );
  HDOAI211DL U1763 ( .A1(n2944), .A2(n2948), .B(n2952), .C(n1601), .Z(n1992)
         );
  HDNAN2D2 U1764 ( .A1(n2725), .A2(instruction[8]), .Z(n2986) );
  HDAOI21M20D2 U1765 ( .A1(n2316), .A2(n2929), .B(n2315), .Z(n2344) );
  HDAND2DL U1766 ( .A1(n1890), .A2(n1599), .Z(n1915) );
  HDINVDL U1767 ( .A(n930), .Z(n2984) );
  HDINVBD2 U1768 ( .A(n2274), .Z(n2468) );
  HDINVD2 U1769 ( .A(n2001), .Z(n1990) );
  HDOAI222DL U1770 ( .A1(n1737), .A2(n2370), .B1(n2934), .B2(n2369), .C1(n1732), .C2(n2368), .Z(o_m_opcode[5]) );
  HDNOR2D2 U1771 ( .A1(n2085), .A2(n2062), .Z(n2906) );
  HDOAI222DL U1772 ( .A1(n1737), .A2(n2097), .B1(n2934), .B2(n2096), .C1(n1732), .C2(n2095), .Z(o_m_opcode[0]) );
  HDNOR4D2 U1773 ( .A1(n2071), .A2(n2114), .A3(n2070), .A4(n2069), .Z(n2159)
         );
  HDNOR2D2 U1774 ( .A1(n2548), .A2(n2592), .Z(n1680) );
  HDINVD4 U1775 ( .A(n1985), .Z(n2242) );
  HDOAI21M20D2 U1776 ( .A1(n2543), .A2(n1846), .B(n2563), .Z(n2554) );
  HDOA211D2 U1777 ( .A1(n2812), .A2(n1845), .B(n1844), .C(n1843), .Z(n2563) );
  HDINVD1 U1778 ( .A(n387), .Z(n2976) );
  HDOR2D4 U1779 ( .A1(instruction[6]), .A2(instruction[5]), .Z(n387) );
  HDOAI21M20DL U1780 ( .A1(n2017), .A2(n2013), .B(n1609), .Z(n2014) );
  HDNOR3D2 U1781 ( .A1(n2624), .A2(n2605), .A3(n2004), .Z(n1679) );
  HDAND4D2 U1782 ( .A1(n1676), .A2(n1997), .A3(n1677), .A4(n1720), .Z(n2004)
         );
  HDNOR2D2 U1783 ( .A1(instruction[11]), .A2(n2978), .Z(n1161) );
  HDNAN2D2 U1784 ( .A1(n2550), .A2(n2005), .Z(n2212) );
  HDOR2D4 U1785 ( .A1(n2242), .A2(n1689), .Z(n2550) );
  HDNAN2D2 U1786 ( .A1(n2161), .A2(n2001), .Z(n2005) );
  HDINVD2 U1787 ( .A(n1689), .Z(n2161) );
  HDNAN3D2 U1788 ( .A1(n1681), .A2(n1682), .A3(n1683), .Z(o_m_futype[2]) );
  HDINVD2 U1789 ( .A(o_m_branch_type[3]), .Z(n1681) );
  HDMUXB2D1 U1790 ( .A0(n1654), .A1(n2947), .SL(n2696), .Z(n1653) );
  HDOR2D4 U1791 ( .A1(n1707), .A2(n1708), .Z(n2927) );
  HDNAN4DL U1792 ( .A1(n2025), .A2(n2525), .A3(n2930), .A4(n2140), .Z(n1870)
         );
  HDOAI211D1 U1793 ( .A1(n2950), .A2(n1689), .B(n2948), .C(n1600), .Z(o_rd[2])
         );
  HDNAN4D1 U1794 ( .A1(n2631), .A2(n2562), .A3(n2588), .A4(n2596), .Z(n2566)
         );
  HDNOR3D1 U1795 ( .A1(n2866), .A2(n2865), .A3(n2864), .Z(n1651) );
  HDOAI211D1 U1796 ( .A1(n2222), .A2(n2377), .B(n2221), .C(n2220), .Z(n2223)
         );
  HDNAN3DL U1797 ( .A1(n2619), .A2(n2216), .A3(n2215), .Z(n2218) );
  HDNOR2D1 U1798 ( .A1(n2597), .A2(n2346), .Z(n2429) );
  HDNOR4D1 U1799 ( .A1(n2454), .A2(n2410), .A3(n2762), .A4(n2409), .Z(n2433)
         );
  HDNOR4D1 U1800 ( .A1(n1821), .A2(n2883), .A3(n1820), .A4(n1877), .Z(n1698)
         );
  HDAOI21M20DL U1801 ( .A1(n2241), .A2(n1812), .B(n2501), .Z(n1813) );
  HDOAI31D1 U1802 ( .A1(n2326), .A2(n2325), .A3(n2324), .B(n2323), .Z(n1629)
         );
  HDNAN2D1 U1803 ( .A1(n2725), .A2(n2685), .Z(n1639) );
  HDNAN4D1 U1804 ( .A1(n2875), .A2(n2874), .A3(n2873), .A4(n2872), .Z(n2877)
         );
  HDNOR3D1 U1805 ( .A1(n2871), .A2(n2870), .A3(n2869), .Z(n2875) );
  HDAOI22D1 U1806 ( .A1(n2348), .A2(n2423), .B1(n2347), .B2(n2597), .Z(n2350)
         );
  HDAOI21D1 U1807 ( .A1(n2982), .A2(n2981), .B(instruction[8]), .Z(n922) );
  HDAOI222D1 U1808 ( .A1(n2296), .A2(n2295), .B1(n2294), .B2(n2293), .C1(n2292), .C2(n2881), .Z(n2297) );
  HDAND2DL U1809 ( .A1(n2186), .A2(n2399), .Z(n2315) );
  HDNAN4DL U1810 ( .A1(n2271), .A2(n2260), .A3(n2259), .A4(n2582), .Z(n2261)
         );
  HDNAN4D1 U1811 ( .A1(n2641), .A2(n2673), .A3(n2767), .A4(n2640), .Z(n2642)
         );
  HDNOR3D1 U1812 ( .A1(n2667), .A2(n2789), .A3(n2666), .Z(n2694) );
  HDAOI211D1 U1813 ( .A1(n2982), .A2(n2981), .B(instruction[8]), .C(
        instruction[7]), .Z(n1094) );
  HDAOI211DL U1814 ( .A1(n2322), .A2(instruction[26]), .B(n2153), .C(n2152), 
        .Z(n2154) );
  HDAOI211D1 U1815 ( .A1(n2778), .A2(n1685), .B(n2667), .C(n2141), .Z(n2142)
         );
  HDINVD1 U1816 ( .A(n1133), .Z(n2109) );
  HDMUX2D1 U1817 ( .A0(n2102), .A1(n2101), .SL(instruction[12]), .Z(n2163) );
  HDAOI211DL U1818 ( .A1(n1701), .A2(n2795), .B(n2773), .C(n425), .Z(n2776) );
  HDNAN3DL U1819 ( .A1(n2820), .A2(n2083), .A3(n2418), .Z(n2084) );
  HDNOR2D1 U1820 ( .A1(n2435), .A2(n1686), .Z(n2280) );
  HDNOR2D1 U1821 ( .A1(n2041), .A2(n2040), .Z(n2043) );
  HDNOR2D1 U1822 ( .A1(n2499), .A2(n2373), .Z(n2044) );
  HDNAN2D1 U1823 ( .A1(n2121), .A2(n2019), .Z(n2191) );
  HDINVD1 U1824 ( .A(n2482), .Z(n2020) );
  HDINVD1 U1825 ( .A(n2789), .Z(n2930) );
  HDNOR2D1 U1826 ( .A1(n2102), .A2(n1947), .Z(n2727) );
  HDNAN2D1 U1827 ( .A1(n2478), .A2(n1599), .Z(n2840) );
  HDNOR2D1 U1828 ( .A1(instruction[17]), .A2(instruction[18]), .Z(n2771) );
  HDINVBD4 U1829 ( .A(instruction[16]), .Z(n2810) );
  HDINVD1 U1830 ( .A(n2282), .Z(n2537) );
  HDINVBD2 U1831 ( .A(n2502), .Z(n2870) );
  HDNAN2D1 U1832 ( .A1(n2676), .A2(n2418), .Z(n2734) );
  HDNAN3D1 U1833 ( .A1(n1888), .A2(instruction[19]), .A3(n2374), .Z(n2732) );
  HDNAN2M1D2 U1834 ( .A1(n2578), .A2(n2501), .Z(n2502) );
  HDNOR2D1 U1835 ( .A1(n1861), .A2(n2578), .Z(n2864) );
  HDAOI21D1 U1836 ( .A1(n2677), .A2(n2495), .B(n1736), .Z(o_m_type[2]) );
  HDNOR2D2 U1837 ( .A1(n2578), .A2(n1831), .Z(n2408) );
  HDNAN2D2 U1838 ( .A1(n2696), .A2(instruction[26]), .Z(n2943) );
  HDNOR2D2 U1839 ( .A1(n2944), .A2(n1990), .Z(n2325) );
  HDNOR2D6 U1840 ( .A1(n1864), .A2(instruction[13]), .Z(n2881) );
  HDNOR2D1 U1841 ( .A1(n1137), .A2(instruction[7]), .Z(n840) );
  HDINVD1 U1842 ( .A(n1702), .Z(n1137) );
  HDNAN2D1 U1843 ( .A1(n2706), .A2(n2705), .Z(n2708) );
  HDNAN2D2 U1844 ( .A1(instruction[11]), .A2(instruction[10]), .Z(n2102) );
  HDNAN2D2 U1845 ( .A1(n2501), .A2(n1731), .Z(n2524) );
  HDNAN2D4 U1846 ( .A1(n1772), .A2(n2812), .Z(n2597) );
  HDNAN2D2 U1847 ( .A1(n2444), .A2(n2811), .Z(n2270) );
  HDNOR2D2 U1848 ( .A1(instruction[27]), .A2(instruction[26]), .Z(n2336) );
  HDAND2D1 U1849 ( .A1(n1823), .A2(n1822), .Z(n2644) );
  HDNAN2D1 U1850 ( .A1(n2493), .A2(n2659), .Z(n2186) );
  HDNAN2D1 U1851 ( .A1(n2500), .A2(n2257), .Z(n1879) );
  HDINVD8 U1852 ( .A(instruction[22]), .Z(n1951) );
  HDOAI31D1 U1853 ( .A1(n1875), .A2(n1732), .A3(n2064), .B(n1872), .Z(
        o_m_ccshift[1]) );
  HDNAN3DL U1854 ( .A1(n2590), .A2(n2589), .A3(n2952), .Z(n2591) );
  HDNOR4D1 U1855 ( .A1(n2276), .A2(n2275), .A3(n591), .A4(n2291), .Z(n2277) );
  HDOAI211D1 U1856 ( .A1(n1879), .A2(instruction[25]), .B(n2422), .C(n2475), 
        .Z(n2252) );
  HDINVDL U1857 ( .A(n2377), .Z(n2235) );
  HDAOI21M20DL U1858 ( .A1(n2658), .A2(n2732), .B(n2384), .Z(n2751) );
  HDNAN2D2 U1859 ( .A1(n2505), .A2(n2812), .Z(n2443) );
  HDAO31DL U1860 ( .A1(n2776), .A2(n2775), .A3(n2774), .B(n1732), .Z(n2780) );
  HDAOI211D1 U1861 ( .A1(n2481), .A2(n2784), .B(n2049), .C(n2048), .Z(n2050)
         );
  HDNOR3D1 U1862 ( .A1(n2282), .A2(instruction[14]), .A3(n2810), .Z(n2540) );
  HDNOR2D2 U1863 ( .A1(instruction[15]), .A2(instruction[16]), .Z(n2310) );
  HDNOR2D2 U1864 ( .A1(n2486), .A2(n2460), .Z(n2437) );
  HDINVD1 U1865 ( .A(n2927), .Z(n2899) );
  HDNAN3D1 U1866 ( .A1(n1777), .A2(instruction[21]), .A3(n1951), .Z(n2459) );
  HDNAN2D2 U1867 ( .A1(n2500), .A2(n1731), .Z(n2475) );
  HDNAN2DL U1868 ( .A1(n2820), .A2(n2819), .Z(n2821) );
  HDAOI22DL U1869 ( .A1(n2294), .A2(n2984), .B1(n2713), .B2(n2182), .Z(n2164)
         );
  HDNAN3DL U1870 ( .A1(n1093), .A2(n2159), .A3(n2312), .Z(n2169) );
  HDNOR2DL U1871 ( .A1(n2738), .A2(n2617), .Z(n2445) );
  HDINVDL U1872 ( .A(n2435), .Z(n2439) );
  HDOAI21DL U1873 ( .A1(n2336), .A2(n2951), .B(n2321), .Z(n1630) );
  HDNOR2M1DL U1874 ( .A1(n1622), .A2(n2766), .Z(n1621) );
  HDNOR2DL U1875 ( .A1(n2889), .A2(n1736), .Z(n2913) );
  HDNOR2D1 U1876 ( .A1(n2579), .A2(n1736), .Z(n1742) );
  HDNAN4DL U1877 ( .A1(n2286), .A2(n2285), .A3(n1619), .A4(n2284), .Z(n2289)
         );
  HDOAI31DL U1878 ( .A1(n2761), .A2(n2649), .A3(n2648), .B(n1599), .Z(n2651)
         );
  HDINVDL U1879 ( .A(n2674), .Z(n2649) );
  HDNAN4D1 U1880 ( .A1(n2657), .A2(n2656), .A3(n2655), .A4(n2654), .Z(n2668)
         );
  HDNOR2D1 U1881 ( .A1(n2939), .A2(n2977), .Z(n2639) );
  HDNAN2DL U1882 ( .A1(n2985), .A2(n679), .Z(n2276) );
  HDOAI22DL U1883 ( .A1(n644), .A2(n2415), .B1(n2110), .B2(n2927), .Z(n2077)
         );
  HDINVDL U1884 ( .A(n2784), .Z(n2902) );
  HDINVD2 U1885 ( .A(n2986), .Z(n2960) );
  HDAOI22DL U1886 ( .A1(instruction[10]), .A2(instruction[12]), .B1(n2675), 
        .B2(instruction[9]), .Z(n2785) );
  HDINVDL U1887 ( .A(n2543), .Z(n1850) );
  HDNAN3D2 U1888 ( .A1(n2295), .A2(instruction[18]), .A3(n2797), .Z(n2055) );
  HDNAN2D2 U1889 ( .A1(n2560), .A2(n2282), .Z(n2295) );
  HDINVD1 U1890 ( .A(n2384), .Z(n2376) );
  HDNAN3D1 U1891 ( .A1(n2767), .A2(n2733), .A3(n2732), .Z(n2735) );
  HDNAN2DL U1892 ( .A1(n2327), .A2(n2377), .Z(n1981) );
  HDNOR3D4 U1893 ( .A1(n1769), .A2(n2486), .A3(n2586), .Z(n2656) );
  HDNOR3D4 U1894 ( .A1(n2085), .A2(instruction[9]), .A3(n2101), .Z(n2481) );
  HDINVD1 U1895 ( .A(n2147), .Z(n1996) );
  HDINVD1 U1896 ( .A(n2589), .Z(n2619) );
  HDINVD2 U1897 ( .A(n2968), .Z(n835) );
  HDINVBD4 U1898 ( .A(instruction[9]), .Z(n1947) );
  HDNAN2DL U1899 ( .A1(instruction[9]), .A2(n1395), .Z(n1741) );
  HDINVBD4 U1900 ( .A(n2189), .Z(n2579) );
  HDNAN2D4 U1901 ( .A1(n2256), .A2(n1888), .Z(n2767) );
  HDNAN3D1 U1902 ( .A1(n1770), .A2(n1777), .A3(n1951), .Z(n2463) );
  HDNAN2D2 U1903 ( .A1(instruction[24]), .A2(instruction[22]), .Z(n1752) );
  HDNOR3D2 U1904 ( .A1(n1878), .A2(n2082), .A3(n2762), .Z(n2827) );
  HDAOI21DL U1905 ( .A1(n2306), .A2(n2202), .B(n1736), .Z(o_m_access_size[1])
         );
  HDAOI31DL U1906 ( .A1(n2564), .A2(n2597), .A3(n2625), .B(n2628), .Z(n2565)
         );
  HDAND2DL U1907 ( .A1(n2957), .A2(instruction[25]), .Z(o_rd[5]) );
  HDAND4DL U1908 ( .A1(n2558), .A2(n2557), .A3(n2597), .A4(n2625), .Z(n2588)
         );
  HDOR4D1 U1909 ( .A1(n2580), .A2(n2579), .A3(n2977), .A4(n2578), .Z(n2581) );
  HDOR2DL U1910 ( .A1(n2435), .A2(n2658), .Z(n2421) );
  HDOAI222DL U1911 ( .A1(n1619), .A2(n2443), .B1(n2380), .B2(n2767), .C1(n2916), .C2(n2983), .Z(n1634) );
  HDOAI211DL U1912 ( .A1(n2394), .A2(n930), .B(n1639), .C(n1640), .Z(n1638) );
  HDAOI21DL U1913 ( .A1(n2189), .A2(n2139), .B(n2021), .Z(n2306) );
  HDNAN2DL U1914 ( .A1(n2960), .A2(n2706), .Z(n1790) );
  HDNAN2DL U1915 ( .A1(n2451), .A2(n2450), .Z(n2452) );
  HDINVDL U1916 ( .A(n2928), .Z(n2783) );
  HDOAI21M20D1 U1917 ( .A1(n2170), .A2(n644), .B(n2158), .Z(n1758) );
  HDNAN2DL U1918 ( .A1(n2616), .A2(n2598), .Z(n2541) );
  HDNOR3DL U1919 ( .A1(n2929), .A2(n441), .A3(n2988), .Z(n2756) );
  HDNAN2D1 U1920 ( .A1(n2417), .A2(n2443), .Z(n2296) );
  HDNAN2DL U1921 ( .A1(n992), .A2(n2468), .Z(n2275) );
  HDNAN3DL U1922 ( .A1(n2873), .A2(n2495), .A3(n2332), .Z(n2454) );
  HDAND2D2 U1923 ( .A1(n2881), .A2(n2465), .Z(n2360) );
  HDNOR3D1 U1924 ( .A1(n2989), .A2(n2086), .A3(n2085), .Z(n2311) );
  HDNAN2DL U1925 ( .A1(n2968), .A2(n2784), .Z(n2895) );
  HDAOI21M20D1 U1926 ( .A1(n1133), .A2(n1231), .B(n2987), .Z(n2069) );
  HDAOI21M20D1 U1927 ( .A1(n1133), .A2(n990), .B(n2927), .Z(n2070) );
  HDAO22D1 U1928 ( .A1(n2723), .A2(n2705), .B1(n2959), .B2(n2465), .Z(n2111)
         );
  HDNAN2D2 U1929 ( .A1(n2061), .A2(n2883), .Z(n2417) );
  HDOR2DL U1930 ( .A1(n2784), .A2(n2973), .Z(n415) );
  HDNAN2DL U1931 ( .A1(n1873), .A2(n2189), .Z(n2331) );
  HDAND3DL U1932 ( .A1(n2382), .A2(n2259), .A3(n2046), .Z(n2130) );
  HDNOR2D2 U1933 ( .A1(n2927), .A2(n2983), .Z(n2964) );
  HDNAN3DL U1934 ( .A1(n2537), .A2(n2536), .A3(n2797), .Z(n2615) );
  HDNOR2DL U1935 ( .A1(n2943), .A2(n1990), .Z(n2006) );
  HDAOI222DL U1936 ( .A1(n2935), .A2(n2972), .B1(n2805), .B2(n2713), .C1(n2973), .C2(n2712), .Z(n2714) );
  HDINVD2 U1937 ( .A(n441), .Z(n2705) );
  HDINVD2 U1938 ( .A(n2973), .Z(n2755) );
  HDINVBD4 U1939 ( .A(instruction[7]), .Z(n2980) );
  HDAND2D1 U1940 ( .A1(n2189), .A2(n1888), .Z(n2510) );
  HDAND2D2 U1941 ( .A1(n2495), .A2(n2493), .Z(n2674) );
  HDINVDL U1942 ( .A(n2486), .Z(n1853) );
  HDINVD1 U1943 ( .A(n2258), .Z(n1753) );
  HDAOI22DL U1944 ( .A1(n2859), .A2(n2620), .B1(n2846), .B2(n2845), .Z(n2621)
         );
  HDOAI211DL U1945 ( .A1(n2619), .A2(instruction[29]), .B(n2618), .C(n1720), 
        .Z(n2846) );
  HDAND3DL U1946 ( .A1(n2701), .A2(n2464), .A3(n2463), .Z(n2474) );
  HDNOR4DL U1947 ( .A1(n2648), .A2(n2739), .A3(n2499), .A4(n2920), .Z(n1782)
         );
  HDINVDL U1948 ( .A(n2554), .Z(n2631) );
  HDNAN2D1 U1949 ( .A1(n2691), .A2(instruction[27]), .Z(n2688) );
  HDNAN4D1 U1950 ( .A1(n2759), .A2(n2654), .A3(n2202), .A4(n2201), .Z(n2204)
         );
  HDNAN2DL U1951 ( .A1(n2986), .A2(n2170), .Z(n2173) );
  HDNAN3DL U1952 ( .A1(n2881), .A2(n2878), .A3(n409), .Z(n2416) );
  HDAOI21M20DL U1953 ( .A1(n1722), .A2(n1736), .B(n1871), .Z(n1826) );
  HDNAN2M1DL U1954 ( .A1(n1229), .A2(n2928), .Z(n470) );
  HDNOR3DL U1955 ( .A1(n1688), .A2(n2948), .A3(n2946), .Z(n1631) );
  HDAOI211DL U1956 ( .A1(n2658), .A2(n2501), .B(n2522), .C(n2500), .Z(n2514)
         );
  HDOAI21DL U1957 ( .A1(n2389), .A2(n388), .B(n885), .Z(n2353) );
  HDNOR3DL U1958 ( .A1(n2679), .A2(n2336), .A3(n2951), .Z(n2337) );
  HDNAN2DL U1959 ( .A1(n2283), .A2(n2810), .Z(n2286) );
  HDOAI21D1 U1960 ( .A1(n2802), .A2(n2795), .B(n2183), .Z(n2103) );
  HDINVDL U1961 ( .A(n2971), .Z(n2075) );
  HDINVD1 U1962 ( .A(n2522), .Z(n2819) );
  HDOAI22DL U1963 ( .A1(n2972), .A2(n2988), .B1(n671), .B2(n2927), .Z(n1660)
         );
  HDNAN3D2 U1964 ( .A1(n2905), .A2(n1685), .A3(n2723), .Z(n1976) );
  HDINVD1 U1965 ( .A(n2845), .Z(n2604) );
  HDNAN2D1 U1966 ( .A1(n2618), .A2(n2522), .Z(n2551) );
  HDNAN2D1 U1967 ( .A1(n1697), .A2(n2952), .Z(n2618) );
  HDOR2DL U1968 ( .A1(n2266), .A2(n2510), .Z(n1802) );
  HDNAN2D4 U1969 ( .A1(n2171), .A2(n2860), .Z(n2603) );
  HDNAN2DL U1970 ( .A1(n2810), .A2(instruction[15]), .Z(n1849) );
  HDNAN3DL U1971 ( .A1(n2482), .A2(n2259), .A3(n2463), .Z(n1666) );
  HDNAN2DL U1972 ( .A1(n2731), .A2(n2730), .Z(n2736) );
  HDNOR2D2 U1973 ( .A1(n2327), .A2(n1706), .Z(n2834) );
  HDNAN2D1 U1974 ( .A1(n2817), .A2(n2738), .Z(n2920) );
  HDINVD2 U1975 ( .A(n2510), .Z(n2738) );
  HDNOR2D2 U1976 ( .A1(n2406), .A2(n2585), .Z(n1751) );
  HDNOR2D2 U1977 ( .A1(n1750), .A2(n2377), .Z(n2585) );
  HDAOI31D2 U1978 ( .A1(n2017), .A2(n2907), .A3(n2767), .B(n1732), .Z(
        o_m_branch_type[3]) );
  HDNOR2D2 U1979 ( .A1(n2003), .A2(n2002), .Z(n2605) );
  HDNAN4D4 U1980 ( .A1(n2546), .A2(n2032), .A3(n2658), .A4(n2619), .Z(n1999)
         );
  HDNOR2D2 U1981 ( .A1(n2944), .A2(n1986), .Z(n2213) );
  HDINVD2 U1982 ( .A(n1544), .Z(n1806) );
  HDNAN2D1 U1983 ( .A1(n1888), .A2(n2258), .Z(n2128) );
  HDAND2D2 U1984 ( .A1(n2019), .A2(n2450), .Z(n2817) );
  HDNAN2D1 U1985 ( .A1(n1823), .A2(n1888), .Z(n2019) );
  HDNOR2D4 U1986 ( .A1(n2327), .A2(n1831), .Z(n2406) );
  HDNAN2D1 U1987 ( .A1(n2374), .A2(instruction[20]), .Z(n2681) );
  HDAND3D2 U1988 ( .A1(n1822), .A2(n2258), .A3(instruction[23]), .Z(n2040) );
  HDNOR2DL U1989 ( .A1(n1860), .A2(n1736), .Z(o_m_access_size[0]) );
  HDNOR3DL U1990 ( .A1(n1878), .A2(n2082), .A3(n2762), .Z(n1699) );
  HDAOI21M20DL U1991 ( .A1(n2694), .A2(n1736), .B(o_m_access_size_6_), .Z(
        n2697) );
  HDNOR2D2 U1992 ( .A1(n1721), .A2(n2855), .Z(n2915) );
  HDOAI21M20DL U1993 ( .A1(n2800), .A2(n2799), .B(n2798), .Z(n2801) );
  HDNAN3DL U1994 ( .A1(n2577), .A2(n2917), .A3(n2657), .Z(n2587) );
  HDNAN2DL U1995 ( .A1(n2785), .A2(n2784), .Z(n2786) );
  HDOAI211DL U1996 ( .A1(n2960), .A2(n2988), .B(n2783), .C(n2987), .Z(n2788)
         );
  HDAOI211DL U1997 ( .A1(n1706), .A2(n2680), .B(n2934), .C(n2679), .Z(n2682)
         );
  HDINVDL U1998 ( .A(n2764), .Z(n2335) );
  HDAND4D1 U1999 ( .A1(n2577), .A2(n1596), .A3(n2376), .A4(n2656), .Z(n1754)
         );
  HDAOI211D1 U2000 ( .A1(n2543), .A2(n2542), .B(n2556), .C(n2541), .Z(n2544)
         );
  HDNAN2DL U2001 ( .A1(n2784), .A2(n2979), .Z(n2744) );
  HDINVBD2 U2002 ( .A(n2360), .Z(n2852) );
  HDOAI31DL U2003 ( .A1(n2660), .A2(n2739), .A3(n2921), .B(n1599), .Z(n2661)
         );
  HDAND4D1 U2004 ( .A1(n2385), .A2(n2699), .A3(n2437), .A4(n2751), .Z(n2388)
         );
  HDOAI21M20DL U2005 ( .A1(n2241), .A2(n2258), .B(n1731), .Z(n2405) );
  HDNAN2DL U2006 ( .A1(n2659), .A2(n2046), .Z(n2748) );
  HDNAN2DL U2007 ( .A1(n2231), .A2(n2948), .Z(n2321) );
  HDNAN2DL U2008 ( .A1(n1802), .A2(n2265), .Z(n2609) );
  HDNOR3D2 U2009 ( .A1(n2119), .A2(n1842), .A3(n1841), .Z(n1843) );
  HDNOR2D1 U2010 ( .A1(n2543), .A2(instruction[15]), .Z(n1838) );
  HDINVD2 U2011 ( .A(instruction[14]), .Z(n2797) );
  HDNAN2DL U2012 ( .A1(n2323), .A2(n1712), .Z(n2690) );
  HDNAN2D2 U2013 ( .A1(n1596), .A2(n2816), .Z(n2871) );
  HDAO211DL U2014 ( .A1(n1609), .A2(n2698), .B(n2497), .C(o_m_flags[3]), .Z(
        o_m_branch_type[2]) );
  HDNOR2D1 U2015 ( .A1(n2817), .A2(n1732), .Z(o_m_flags[3]) );
  HDNAN3D2 U2016 ( .A1(n1751), .A2(n2472), .A3(n2459), .Z(n1769) );
  HDAOI211D2 U2017 ( .A1(n2009), .A2(o_rs2_1_), .B(n2324), .C(n2008), .Z(n2570) );
  HDNAN2M1DL U2018 ( .A1(instruction[29]), .A2(n1995), .Z(n1678) );
  HDINVBD4 U2019 ( .A(instruction[6]), .Z(n2981) );
  HDINVD2 U2020 ( .A(n633), .Z(n2972) );
  HDNOR2D2 U2021 ( .A1(n2102), .A2(instruction[9]), .Z(n2925) );
  HDNAN2D2 U2022 ( .A1(n2973), .A2(n2980), .Z(n633) );
  HDINVD1 U2023 ( .A(n2767), .Z(n2356) );
  HDINVD1 U2024 ( .A(n2270), .Z(n1772) );
  HDNAN3D2 U2025 ( .A1(n2701), .A2(n2700), .A3(n1611), .Z(n2880) );
  HDAND2D1 U2026 ( .A1(n1596), .A2(n2699), .Z(n1611) );
  HDNOR4D2 U2027 ( .A1(n2462), .A2(n2461), .A3(n2460), .A4(n2644), .Z(n2701)
         );
  HDNOR2D2 U2028 ( .A1(n2499), .A2(n2406), .Z(n2483) );
  HDNOR2D1 U2029 ( .A1(n1812), .A2(n1688), .Z(n2082) );
  HDINVD2 U2030 ( .A(n2501), .Z(n2198) );
  HDNAN3D1 U2031 ( .A1(n2963), .A2(n400), .A3(n2851), .Z(n2856) );
  HDINVDL U2032 ( .A(n2938), .Z(n2807) );
  HDNAN2D1 U2033 ( .A1(n2801), .A2(n1735), .Z(n2814) );
  HDNOR2DL U2034 ( .A1(n2633), .A2(n2632), .Z(n2635) );
  HDINVD1 U2035 ( .A(n2489), .Z(n2487) );
  HDNAN4DL U2036 ( .A1(n2375), .A2(n2951), .A3(n2948), .A4(n2379), .Z(n2207)
         );
  HDNOR2DL U2037 ( .A1(n2282), .A2(instruction[16]), .Z(n2174) );
  HDNOR2DL U2038 ( .A1(n2162), .A2(n2161), .Z(n2165) );
  HDAOI31D1 U2039 ( .A1(n2319), .A2(n2639), .A3(n2389), .B(n1636), .Z(n1635)
         );
  HDINVDL U2040 ( .A(n2932), .Z(n2512) );
  HDNAN4D1 U2041 ( .A1(n2908), .A2(n2956), .A3(n2907), .A4(n2916), .Z(n2909)
         );
  HDOAI21M20D1 U2042 ( .A1(n1797), .A2(n2705), .B(n1758), .Z(n2897) );
  HDAOI21M20D1 U2043 ( .A1(n1920), .A2(n1915), .B(n2978), .Z(n1916) );
  HDNOR2D2 U2044 ( .A1(n2929), .A2(n2987), .Z(n2355) );
  HDAOI22D1 U2045 ( .A1(n2639), .A2(n2354), .B1(n2800), .B2(n2353), .Z(n2358)
         );
  HDNAN2DL U2046 ( .A1(n2614), .A2(n2538), .Z(n2539) );
  HDNAN3DL U2047 ( .A1(n1965), .A2(n1964), .A3(n1957), .Z(o_m_imm[24]) );
  HDNAN3DL U2048 ( .A1(n1965), .A2(n1964), .A3(n1956), .Z(o_m_imm[23]) );
  HDNAN3DL U2049 ( .A1(n1716), .A2(n1964), .A3(n1958), .Z(o_m_imm[25]) );
  HDNAN3DL U2050 ( .A1(n1716), .A2(n1964), .A3(n1960), .Z(o_m_imm[27]) );
  HDNAN3DL U2051 ( .A1(n1716), .A2(n1964), .A3(n1959), .Z(o_m_imm[26]) );
  HDOAI21DL U2052 ( .A1(n2981), .A2(n834), .B(n2313), .Z(n2292) );
  HDAOI22DL U2053 ( .A1(n2447), .A2(n2289), .B1(n2288), .B2(n2287), .Z(n2298)
         );
  HDOAI21DL U2054 ( .A1(n2800), .A2(n2795), .B(n1609), .Z(n2652) );
  HDOAI21M20D1 U2055 ( .A1(n1922), .A2(n1921), .B(n1599), .Z(n1723) );
  HDAOI22DL U2056 ( .A1(n2146), .A2(n2145), .B1(n2144), .B2(n2492), .Z(n2208)
         );
  HDNAN4D1 U2057 ( .A1(n2129), .A2(n2309), .A3(n2482), .A4(n2128), .Z(n2342)
         );
  HDAOI21DL U2058 ( .A1(n2124), .A2(n2811), .B(instruction[15]), .Z(n2127) );
  HDNOR3D1 U2059 ( .A1(n2726), .A2(n591), .A3(n2971), .Z(n2965) );
  HDINVBD4 U2060 ( .A(n2800), .Z(n2901) );
  HDINVDL U2061 ( .A(n2266), .Z(n2107) );
  HDNAN2DL U2062 ( .A1(n1731), .A2(n2189), .Z(n2140) );
  HDNAN3D1 U2063 ( .A1(n2641), .A2(n2819), .A3(n2271), .Z(n1862) );
  HDNAN2DL U2064 ( .A1(n1731), .A2(n1865), .Z(n2046) );
  HDNOR4D1 U2065 ( .A1(n1821), .A2(n2883), .A3(n1820), .A4(n1877), .Z(n1665)
         );
  HDAOI21DL U2066 ( .A1(n2380), .A2(n1981), .B(n2323), .Z(n2016) );
  HDNAN2D2 U2067 ( .A1(n2543), .A2(n2811), .Z(n2560) );
  HDOAI21D1 U2068 ( .A1(n1838), .A2(n1848), .B(n2270), .Z(n1839) );
  HDNAN2D2 U2069 ( .A1(n2511), .A2(n2508), .Z(n1912) );
  HDNOR3D2 U2070 ( .A1(n1885), .A2(n1884), .A3(n1883), .Z(n2763) );
  HDAND3D1 U2071 ( .A1(n2382), .A2(n2475), .A3(n2450), .Z(n1880) );
  HDNAN3D2 U2072 ( .A1(n2731), .A2(n2730), .A3(n1771), .Z(n2862) );
  HDNOR2D2 U2073 ( .A1(n2266), .A2(n1819), .Z(n2508) );
  HDNAN2D1 U2074 ( .A1(n2654), .A2(n2502), .Z(n2503) );
  HDINVD1 U2075 ( .A(n2578), .Z(n2375) );
  HDINVD2 U2076 ( .A(n1865), .Z(n1835) );
  HDNAN3DL U2077 ( .A1(n1749), .A2(n1748), .A3(instruction[21]), .Z(n1750) );
  HDNAN2D2 U2078 ( .A1(n2515), .A2(n2845), .Z(n2017) );
  HDAO31D1 U2079 ( .A1(n2246), .A2(n2233), .A3(n2029), .B(instruction[29]), 
        .Z(n1730) );
  HDINVDL U2080 ( .A(n1701), .Z(n2911) );
  HDNOR3D2 U2081 ( .A1(n1988), .A2(n1994), .A3(n1987), .Z(n2546) );
  HDNAN3DL U2082 ( .A1(n2233), .A2(n2007), .A3(n2245), .Z(n1727) );
  HDNOR2D2 U2083 ( .A1(n2948), .A2(instruction[28]), .Z(n1985) );
  HDNOR2D2 U2084 ( .A1(n2880), .A2(n2749), .Z(n2769) );
  HDNAN2D4 U2085 ( .A1(n1777), .A2(instruction[22]), .Z(n2327) );
  HDNAN2D2 U2086 ( .A1(instruction[21]), .A2(instruction[19]), .Z(n1743) );
  HDNOR2D2 U2087 ( .A1(n2198), .A2(n1687), .Z(n2049) );
  HDBUFD4 U2088 ( .A(n2338), .Z(n1687) );
  HDAOI21M20DL U2089 ( .A1(n2011), .A2(n2128), .B(n2356), .Z(n1980) );
  HDAND3DL U2090 ( .A1(n2563), .A2(n2562), .A3(n2627), .Z(n2564) );
  HDNAN4DL U2091 ( .A1(n2699), .A2(n2490), .A3(n2483), .A4(n2482), .Z(n2484)
         );
  HDNOR4DL U2092 ( .A1(n2175), .A2(n2543), .A3(n2559), .A4(n2174), .Z(n2180)
         );
  HDNAN2D1 U2093 ( .A1(n2841), .A2(n2840), .Z(o_rd2[2]) );
  HDAOI22D1 U2094 ( .A1(n2849), .A2(N5186), .B1(n2839), .B2(n1609), .Z(n2841)
         );
  HDNAN4D1 U2095 ( .A1(n2603), .A2(n2472), .A3(n2628), .A4(n2653), .Z(n1856)
         );
  HDAO211D1 U2096 ( .A1(n2865), .A2(n2744), .B(n2933), .C(n2743), .Z(n2790) );
  HDAND3D1 U2097 ( .A1(n2887), .A2(n2916), .A3(n2907), .Z(n1618) );
  HDAOI21D1 U2098 ( .A1(n2865), .A2(n2979), .B(n2360), .Z(n2363) );
  HDOAI31D1 U2099 ( .A1(n2799), .A2(n2713), .A3(n2319), .B(n2712), .Z(n2184)
         );
  HDOAI211D1 U2100 ( .A1(n2183), .A2(n2182), .B(n2725), .C(n2805), .Z(n2185)
         );
  HDAND3DL U2101 ( .A1(n2483), .A2(n2482), .A3(n2264), .Z(n1616) );
  HDAOI21DL U2102 ( .A1(n2246), .A2(n2245), .B(n1687), .Z(n2247) );
  HDOAI22M10DL U2103 ( .A1(n2668), .A2(n1701), .B1(n2659), .B2(n2658), .Z(
        n2660) );
  HDAOI22D1 U2104 ( .A1(n1609), .A2(n2664), .B1(n2687), .B2(n2781), .Z(n2662)
         );
  HDAND2DL U2105 ( .A1(n2650), .A2(n1599), .Z(o_rd_type[3]) );
  HDAOI21M20D2 U2106 ( .A1(n2647), .A2(n1732), .B(n2646), .Z(n2670) );
  HDNOR2D2 U2107 ( .A1(n1928), .A2(n1877), .Z(n1898) );
  HDNOR3D4 U2108 ( .A1(n1591), .A2(n1943), .A3(n1728), .Z(n1949) );
  HDNAN4D1 U2109 ( .A1(n2131), .A2(n2130), .A3(n399), .A4(n2604), .Z(n2132) );
  HDNOR3D1 U2110 ( .A1(n2342), .A2(n2384), .A3(n2634), .Z(n2131) );
  HDNOR3D1 U2111 ( .A1(n2311), .A2(n2087), .A3(n2590), .Z(n2090) );
  HDNOR4D1 U2112 ( .A1(n2084), .A2(n2778), .A3(n2859), .A4(n2864), .Z(n2091)
         );
  HDOAI21M20D1 U2113 ( .A1(n2100), .A2(n1811), .B(n2800), .Z(n2359) );
  HDOAI22D1 U2114 ( .A1(n2976), .A2(n2060), .B1(n2059), .B2(n2058), .Z(n2061)
         );
  HDNAN3DL U2115 ( .A1(n2055), .A2(n2054), .A3(n2053), .Z(n2056) );
  HDINVDL U2116 ( .A(n2418), .Z(n2027) );
  HDNAN4D1 U2117 ( .A1(n2022), .A2(n2502), .A3(n2655), .A4(n2422), .Z(n2138)
         );
  HDNOR4D1 U2118 ( .A1(n2021), .A2(n2789), .A3(n2020), .A4(n2191), .Z(n2022)
         );
  HDAND2D2 U2119 ( .A1(n2784), .A2(instruction[7]), .Z(n2725) );
  HDAOI211D1 U2120 ( .A1(n674), .A2(n2723), .B(n2722), .C(n2721), .Z(n1661) );
  HDNAN2D1 U2121 ( .A1(n2113), .A2(instruction[7]), .Z(n2720) );
  HDNOR3D2 U2122 ( .A1(n1976), .A2(n2597), .A3(n2423), .Z(n2241) );
  HDNOR2D2 U2123 ( .A1(n2861), .A2(n2611), .Z(n2530) );
  HDINVD2 U2124 ( .A(n399), .Z(n2611) );
  HDINVD2 U2125 ( .A(n2551), .Z(n2590) );
  HDNAN2D2 U2126 ( .A1(n2545), .A2(n2602), .Z(n2171) );
  HDNOR2D2 U2127 ( .A1(n1852), .A2(n2561), .Z(n2602) );
  HDNOR2D2 U2128 ( .A1(n2554), .A2(n1851), .Z(n2633) );
  HDNOR2D2 U2129 ( .A1(n2811), .A2(instruction[14]), .Z(n1846) );
  HDNAN2D2 U2130 ( .A1(n2811), .A2(instruction[15]), .Z(n2282) );
  HDOA21M10D2 U2131 ( .A2(n1914), .A1(n1733), .B(n1729), .Z(n1726) );
  HDNOR2D2 U2132 ( .A1(n1878), .A2(n2870), .Z(n2764) );
  HDNOR2D2 U2133 ( .A1(n1942), .A2(n1941), .Z(n1974) );
  HDNOR2D2 U2134 ( .A1(n1929), .A2(n2399), .Z(n1941) );
  HDNAN2D2 U2135 ( .A1(n1667), .A2(n1599), .Z(n1929) );
  HDNOR4D2 U2136 ( .A1(n2736), .A2(n2749), .A3(n2735), .A4(n2734), .Z(n2931)
         );
  HDNAN3D1 U2137 ( .A1(n2264), .A2(n2309), .A3(n2327), .Z(n1768) );
  HDINVD2 U2138 ( .A(n2586), .Z(n2264) );
  HDNAN3D2 U2139 ( .A1(n2656), .A2(n2654), .A3(n2673), .Z(n2648) );
  HDNAN2D4 U2140 ( .A1(n2784), .A2(n2980), .Z(n388) );
  HDNOR2D2 U2141 ( .A1(n2951), .A2(instruction[27]), .Z(n2001) );
  HDINVBD2 U2142 ( .A(n2739), .Z(n1864) );
  HDNOR2D2 U2143 ( .A1(n387), .A2(n2979), .Z(n2113) );
  HDNAN2D2 U2144 ( .A1(n2925), .A2(n2399), .Z(n2988) );
  HDOAI22DL U2145 ( .A1(n2018), .A2(n2501), .B1(n2145), .B2(n1777), .Z(n1860)
         );
  HDNOR2D2 U2146 ( .A1(n2522), .A2(n2373), .Z(n2889) );
  HDINVBD2 U2147 ( .A(n1823), .Z(n1861) );
  HDNOR2D4 U2148 ( .A1(n1774), .A2(n1746), .Z(n1865) );
  HDNAN2D2 U2149 ( .A1(n1873), .A2(n2258), .Z(n2464) );
  HDNAN2D2 U2150 ( .A1(n1873), .A2(n2501), .Z(n2482) );
  HDNAN4D1 U2151 ( .A1(n2458), .A2(n2483), .A3(n2863), .A4(n2817), .Z(n2462)
         );
  HDNOR2D6 U2152 ( .A1(n1740), .A2(n1951), .Z(n1888) );
  HDNOR2D2 U2153 ( .A1(n2384), .A2(n2186), .Z(n2863) );
  HDNAN3D2 U2154 ( .A1(n1832), .A2(n2435), .A3(n2361), .Z(n2762) );
  HDNOR2D2 U2155 ( .A1(n2578), .A2(n1713), .Z(n2486) );
  HDINVD2 U2156 ( .A(n1712), .Z(n1713) );
  HDNAN2D8 U2157 ( .A1(n1745), .A2(instruction[22]), .Z(n2578) );
  HDNAN2D2 U2158 ( .A1(n2254), .A2(n2330), .Z(n1878) );
  HDNOR3D2 U2159 ( .A1(n2049), .A2(n2042), .A3(n2040), .Z(n2254) );
  HDNAN2D2 U2160 ( .A1(n1745), .A2(n1951), .Z(n2338) );
  HDINVBD4 U2161 ( .A(instruction[23]), .Z(n1739) );
  HDAOI31DL U2162 ( .A1(n2674), .A2(n2938), .A3(n2673), .B(n1736), .Z(
        o_rs3_type[2]) );
  HDNAN3DL U2163 ( .A1(n1873), .A2(instruction[21]), .A3(n2941), .Z(n1874) );
  HDAOI21M20DL U2164 ( .A1(n2761), .A2(n1696), .B(n1737), .Z(o_m_flags[5]) );
  HDAOI21M20D1 U2165 ( .A1(n1784), .A2(n2934), .B(n1783), .Z(n378) );
  HDAOI21DL U2166 ( .A1(n2323), .A2(n2678), .B(n2322), .Z(n1784) );
  HDAOI22D1 U2167 ( .A1(n2849), .A2(N5187), .B1(n2842), .B2(n1609), .Z(n2844)
         );
  HDNAN3DL U2168 ( .A1(n2590), .A2(n1701), .A3(n2948), .Z(n2568) );
  HDNAN4DL U2169 ( .A1(n1876), .A2(n2863), .A3(n2702), .A4(n2601), .Z(n1830)
         );
  HDAOI22D1 U2170 ( .A1(n2849), .A2(n2696), .B1(n2831), .B2(n1609), .Z(n2833)
         );
  HDOAI21M20D1 U2171 ( .A1(n1718), .A2(n2845), .B(n2623), .Z(n2848) );
  HDNAN4DL U2172 ( .A1(n2328), .A2(n2674), .A3(n2264), .A4(n2464), .Z(n2203)
         );
  HDOAI211DL U2173 ( .A1(n2199), .A2(n2198), .B(n2346), .C(n2332), .Z(n2205)
         );
  HDOAI222D1 U2174 ( .A1(n2166), .A2(n2318), .B1(n2767), .B2(n2165), .C1(n2901), .C2(n2164), .Z(n2167) );
  HDNAN3DL U2175 ( .A1(n2699), .A2(n2863), .A3(n2437), .Z(n2438) );
  HDAND3D1 U2176 ( .A1(n2456), .A2(n2518), .A3(n2828), .Z(n1612) );
  HDOAI222D1 U2177 ( .A1(n2916), .A2(n2979), .B1(n2064), .B2(n1875), .C1(n2980), .C2(n2393), .Z(n1816) );
  HDOAI22DL U2178 ( .A1(n2939), .A2(n387), .B1(n2798), .B2(n1806), .Z(n1817)
         );
  HDOAI211D1 U2179 ( .A1(n1805), .A2(n1864), .B(n1804), .C(n1803), .Z(n1818)
         );
  HDNAN2DL U2180 ( .A1(n1802), .A2(n1715), .Z(n1803) );
  HDINVDL U2181 ( .A(n1910), .Z(n1804) );
  HDAOI211D1 U2182 ( .A1(n2800), .A2(n1638), .B(n2311), .C(n919), .Z(n1637) );
  HDNOR4D4 U2183 ( .A1(n1608), .A2(n1942), .A3(n1941), .A4(n1728), .Z(n1938)
         );
  HDOAI21D1 U2184 ( .A1(n424), .A2(n425), .B(n1609), .Z(n2715) );
  HDOAI21D1 U2185 ( .A1(n1856), .A2(n1855), .B(n1609), .Z(n1857) );
  HDNAN4DL U2186 ( .A1(n2529), .A2(n2530), .A3(n2730), .A4(n1854), .Z(n1855)
         );
  HDINVD1 U2187 ( .A(n2840), .Z(n1837) );
  HDNAN2DL U2188 ( .A1(n2923), .A2(n2789), .Z(n2792) );
  HDAOI21D1 U2189 ( .A1(n2890), .A2(n1609), .B(n2913), .Z(n2891) );
  HDOAI21M20DL U2190 ( .A1(n1893), .A2(o_rs2_1_), .B(n1905), .Z(o_m_imm[1]) );
  HDAOI211D2 U2191 ( .A1(n1609), .A2(n1891), .B(n1913), .C(n1908), .Z(n1905)
         );
  HDNAN2DL U2192 ( .A1(n2894), .A2(n1701), .Z(n2908) );
  HDAOI22D1 U2193 ( .A1(n2356), .A2(n2380), .B1(n2355), .B2(n874), .Z(n2357)
         );
  HDNAN2D1 U2194 ( .A1(n2548), .A2(n2845), .Z(n2549) );
  HDOAI21M20D1 U2195 ( .A1(n1609), .A2(n2356), .B(n1907), .Z(n1900) );
  HDAOI21M20D2 U2196 ( .A1(n1898), .A2(n1732), .B(n1915), .Z(n1907) );
  HDAOI211D2 U2197 ( .A1(n1609), .A2(n1891), .B(n1913), .C(n1908), .Z(n1709)
         );
  HDOAI22DL U2198 ( .A1(n1701), .A2(n2798), .B1(n2852), .B2(n2755), .Z(n2757)
         );
  HDOAI21DL U2199 ( .A1(instruction[14]), .A2(n2282), .B(n2281), .Z(n2283) );
  HDNAN4DL U2200 ( .A1(n2255), .A2(n2254), .A3(n2817), .A4(n2253), .Z(n2262)
         );
  HDAOI21DL U2201 ( .A1(n2244), .A2(n2550), .B(n2243), .Z(n2248) );
  HDOAI31D1 U2202 ( .A1(n2242), .A2(n2578), .A3(n2946), .B(n2405), .Z(n2249)
         );
  HDNAN4D1 U2203 ( .A1(n2670), .A2(n2662), .A3(n2661), .A4(n2695), .Z(
        o_rs3_type[0]) );
  HDNAN4D1 U2204 ( .A1(n2670), .A2(n2652), .A3(n2651), .A4(n2954), .Z(
        o_rs3_valid) );
  HDAND4D1 U2205 ( .A1(n2305), .A2(n2817), .A3(n2819), .A4(n2471), .Z(n2385)
         );
  HDAOI211D2 U2206 ( .A1(n1609), .A2(n1891), .B(n1913), .C(n1908), .Z(n1710)
         );
  HDOAI21DL U2207 ( .A1(n2148), .A2(n2147), .B(n2492), .Z(n2149) );
  HDAOI211D1 U2208 ( .A1(n2865), .A2(n2276), .B(n2106), .C(n2105), .Z(n2123)
         );
  HDNOR2D2 U2209 ( .A1(n388), .A2(instruction[8]), .Z(n2971) );
  HDAOI211D1 U2210 ( .A1(n2771), .A2(n2797), .B(n2057), .C(n2056), .Z(n2081)
         );
  HDNAN4D1 U2211 ( .A1(n2024), .A2(n2130), .A3(n2023), .A4(n2475), .Z(n2028)
         );
  HDNOR3D1 U2212 ( .A1(n2377), .A2(n2934), .A3(n2374), .Z(n1970) );
  HDNOR2D4 U2213 ( .A1(n2059), .A2(n2939), .Z(n2800) );
  HDOAI21D1 U2214 ( .A1(n1655), .A2(n1737), .B(n2934), .Z(n1664) );
  HDNOR2D1 U2215 ( .A1(o_m_flags[3]), .A2(n2770), .Z(n2015) );
  HDNAN2D1 U2216 ( .A1(n2532), .A2(n1609), .Z(n2534) );
  HDNAN3D1 U2217 ( .A1(n2241), .A2(n2323), .A3(n2500), .Z(n2305) );
  HDOAI21M20D1 U2218 ( .A1(n1850), .A2(n1849), .B(n2542), .Z(n2625) );
  HDAOI21D1 U2219 ( .A1(n1921), .A2(n1922), .B(n250), .Z(n1608) );
  HDNAN2M1DL U2220 ( .A1(n1920), .A2(n1929), .Z(n1923) );
  HDINVBD4 U2221 ( .A(n1726), .Z(n1728) );
  HDNAN2D2 U2222 ( .A1(n1974), .A2(n1673), .Z(n1966) );
  HDINVBD4 U2223 ( .A(n2939), .Z(n2883) );
  HDNAN4D1 U2224 ( .A1(n1880), .A2(n2674), .A3(n2655), .A4(n2676), .Z(n1885)
         );
  HDAOI211D1 U2225 ( .A1(n2510), .A2(n1715), .B(n2795), .C(n2737), .Z(n2932)
         );
  HDAOI31D1 U2226 ( .A1(n2867), .A2(n2525), .A3(n2524), .B(n1736), .Z(n2526)
         );
  HDNAN3D1 U2227 ( .A1(n2521), .A2(n2520), .A3(n2582), .Z(n2869) );
  HDINVD2 U2228 ( .A(n2408), .Z(n2654) );
  HDAOI22D1 U2229 ( .A1(n2492), .A2(n2941), .B1(n1684), .B2(n1609), .Z(n1682)
         );
  HDNOR2D2 U2230 ( .A1(n2939), .A2(n2935), .Z(n2865) );
  HDNAN3DL U2231 ( .A1(n2465), .A2(n2979), .A3(n387), .Z(n2466) );
  HDNOR2D4 U2232 ( .A1(n1705), .A2(instruction[5]), .Z(n2784) );
  HDINVD2 U2233 ( .A(instruction[6]), .Z(n1705) );
  HDNAN2DL U2234 ( .A1(n2007), .A2(n1715), .Z(n2008) );
  HDOA211D1 U2235 ( .A1(n2911), .A2(n1689), .B(n2658), .C(n1730), .Z(n2592) );
  HDNOR2D2 U2236 ( .A1(n2696), .A2(instruction[26]), .Z(n2231) );
  HDNAN2M1D4 U2237 ( .A1(n2243), .A2(n2018), .Z(n2939) );
  HDNAN2D2 U2238 ( .A1(n2935), .A2(n2977), .Z(n2059) );
  HDNAN2D4 U2239 ( .A1(n2969), .A2(n2399), .Z(n2987) );
  HDNOR2D2 U2240 ( .A1(n1806), .A2(instruction[9]), .Z(n2969) );
  HDNOR3D1 U2241 ( .A1(n2478), .A2(n2348), .A3(n2042), .Z(n1778) );
  HDNOR2D2 U2242 ( .A1(n1753), .A2(n1869), .Z(n2373) );
  HDNOR3D1 U2243 ( .A1(n2892), .A2(n2650), .A3(n2409), .Z(n1776) );
  HDNAN2D1 U2244 ( .A1(n2655), .A2(n2450), .Z(n2409) );
  HDNOR2D2 U2245 ( .A1(n1812), .A2(n2243), .Z(n2650) );
  HDINVBD4 U2246 ( .A(n2494), .Z(n2511) );
  HDNAN2D2 U2247 ( .A1(n2938), .A2(n2418), .Z(n2494) );
  HDNOR2D2 U2248 ( .A1(n2789), .A2(n2739), .Z(n2938) );
  HDNAN3D2 U2249 ( .A1(n2500), .A2(n1748), .A3(n1951), .Z(n2309) );
  HDOA21M20D2 U2250 ( .A1(instruction[6]), .A2(instruction[5]), .B(n2607), .Z(
        n2861) );
  HDNAN2D2 U2251 ( .A1(n2789), .A2(n1422), .Z(n2085) );
  HDINVD2 U2252 ( .A(n2505), .Z(n2640) );
  HDAND2D2 U2253 ( .A1(n1865), .A2(n2323), .Z(n2795) );
  HDOR2D2 U2254 ( .A1(n2845), .A2(n2522), .Z(n2749) );
  HDAND2D4 U2255 ( .A1(n2322), .A2(n2258), .Z(n2522) );
  HDINVBD2 U2256 ( .A(n2243), .Z(n2322) );
  HDNOR2D4 U2257 ( .A1(n2243), .A2(n1868), .Z(n2845) );
  HDNAN2D2 U2258 ( .A1(n1701), .A2(n2336), .Z(n2509) );
  HDNOR2D2 U2259 ( .A1(instruction[28]), .A2(instruction[29]), .Z(n2893) );
  HDNAN2D2 U2260 ( .A1(n2475), .A2(n2673), .Z(n2384) );
  HDBUFD8 U2261 ( .A(n2240), .Z(n1731) );
  HDNOR3D2 U2262 ( .A1(n1748), .A2(instruction[23]), .A3(instruction[22]), .Z(
        n2240) );
  HDINVBD4 U2263 ( .A(instruction[24]), .Z(n1748) );
  HDNOR3D4 U2264 ( .A1(n2374), .A2(instruction[19]), .A3(instruction[20]), .Z(
        n1823) );
  HDNOR2D4 U2265 ( .A1(n2681), .A2(n1746), .Z(n2500) );
  HDNOR2D2 U2266 ( .A1(n1739), .A2(instruction[24]), .Z(n1745) );
  HDINVBD4 U2267 ( .A(instruction[19]), .Z(n1746) );
  HDNAN2D1 U2268 ( .A1(n1600), .A2(n2951), .Z(o_rd[3]) );
  HDOAI21D1 U2269 ( .A1(n1875), .A2(n1931), .B(n1874), .Z(o_m_ccshift[2]) );
  HDOAI211D1 U2270 ( .A1(n1980), .A2(n1732), .B(n1979), .C(n1978), .Z(
        o_m_branch_type[0]) );
  HDNAN3D1 U2271 ( .A1(n2339), .A2(n2235), .A3(n2941), .Z(n1978) );
  HDNOR2D1 U2272 ( .A1(n2496), .A2(o_m_flags[3]), .Z(n1979) );
  HDOAI21D1 U2273 ( .A1(n2830), .A2(n2828), .B(n2829), .Z(o_rd2_type[0]) );
  HDOAI21M10D1 U2274 ( .A1(n1699), .A2(n2826), .B(n1609), .Z(n2829) );
  HDNOR3D1 U2275 ( .A1(N5188), .A2(N5187), .A3(N5189), .Z(n2830) );
  HDNAN3D1 U2276 ( .A1(n2846), .A2(n2845), .A3(n1734), .Z(n2847) );
  HDINVD1 U2277 ( .A(n2947), .Z(n2950) );
  HDNOR2D1 U2278 ( .A1(n2621), .A2(n1732), .Z(o_rs4[4]) );
  HDNAN3D1 U2279 ( .A1(n2616), .A2(n2615), .A3(n2614), .Z(n2620) );
  HDINVD1 U2280 ( .A(n1871), .Z(n1872) );
  HDNOR4D1 U2281 ( .A1(n2861), .A2(n2823), .A3(n2822), .A4(n2821), .Z(n2825)
         );
  HDOAI211D1 U2282 ( .A1(n2838), .A2(n1732), .B(n2843), .C(n2837), .Z(o_rd2[1]) );
  HDNAN2D1 U2283 ( .A1(n2849), .A2(N5185), .Z(n2837) );
  HDNOR2D1 U2284 ( .A1(n2835), .A2(n2834), .Z(n2838) );
  HDOAI21D1 U2285 ( .A1(n2697), .A2(n2696), .B(n2695), .Z(o_rs3[5]) );
  HDAND2D1 U2286 ( .A1(n2734), .A2(n1599), .Z(o_m_access_size_6_) );
  HDOAI211D1 U2287 ( .A1(n2915), .A2(n1732), .B(n2955), .C(n2914), .Z(
        o_rd_type[2]) );
  HDINVD1 U2288 ( .A(n2913), .Z(n2914) );
  HDNAN4D1 U2289 ( .A1(n2474), .A2(n2473), .A3(n2472), .A4(n2471), .Z(n2479)
         );
  HDINVD1 U2290 ( .A(n1732), .Z(n1734) );
  HDOR3D1 U2291 ( .A1(n2663), .A2(n2797), .A3(n1732), .Z(n379) );
  HDNOR3D1 U2292 ( .A1(n1782), .A2(n2696), .A3(n1736), .Z(n1783) );
  HDNAN2D1 U2293 ( .A1(n2844), .A2(n2843), .Z(o_rd2[3]) );
  HDOAI22D1 U2294 ( .A1(n2946), .A2(n2814), .B1(n2813), .B2(n2809), .Z(
        o_rs1[1]) );
  HDOAI22D1 U2295 ( .A1(n2951), .A2(n2814), .B1(n2813), .B2(n2811), .Z(
        o_rs1[3]) );
  HDOAI22D1 U2296 ( .A1(n2952), .A2(n2814), .B1(n2813), .B2(n2812), .Z(
        o_rs1[4]) );
  HDAOI22D1 U2297 ( .A1(n1732), .A2(n2576), .B1(n2575), .B2(n2574), .Z(
        o_rs4[1]) );
  HDNOR3D1 U2298 ( .A1(n2835), .A2(n2573), .A3(n2572), .Z(n2574) );
  HDINVD1 U2299 ( .A(n2571), .Z(n2573) );
  HDOAI211D1 U2300 ( .A1(n2570), .A2(n2604), .B(n2569), .C(n2568), .Z(n2835)
         );
  HDAOI211D1 U2301 ( .A1(n2567), .A2(n2566), .B(n2565), .C(o_m_flags[2]), .Z(
        n2575) );
  HDNOR2D1 U2302 ( .A1(n2747), .A2(n2746), .Z(o_rs2[0]) );
  HDNOR4D1 U2303 ( .A1(n2745), .A2(n1732), .A3(n2808), .A4(n2790), .Z(n2747)
         );
  HDOAI211D1 U2304 ( .A1(n2729), .A2(n2929), .B(n2798), .C(n2728), .Z(n2745)
         );
  HDNAN2M1D1 U2305 ( .A1(n1647), .A2(n1648), .Z(o_rd_valid) );
  HDNAN2M1D1 U2306 ( .A1(n1732), .A2(n1649), .Z(n1648) );
  HDNAN4D1 U2307 ( .A1(n2915), .A2(n2863), .A3(n1650), .A4(n1651), .Z(n1649)
         );
  HDNOR2M1D1 U2308 ( .A1(n2879), .A2(n2862), .Z(n1650) );
  HDAOI21M10D1 U2309 ( .A1(n2886), .A2(n2854), .B(n2853), .Z(n2855) );
  HDAO21D1 U2310 ( .A1(n2881), .A2(n2857), .B(n2856), .Z(n1721) );
  HDOAI211D1 U2311 ( .A1(n2850), .A2(n2927), .B(n587), .C(n2926), .Z(n2857) );
  HDINVD1 U2312 ( .A(n2964), .Z(n2926) );
  HDAO21D1 U2313 ( .A1(n2974), .A2(n2158), .B(n2897), .Z(n594) );
  HDNOR2D1 U2314 ( .A1(n2974), .A2(n590), .Z(n2850) );
  HDOAI211D1 U2315 ( .A1(n2867), .A2(n1736), .B(n1600), .C(n2868), .Z(n1647)
         );
  HDOAI21D1 U2316 ( .A1(n1897), .A2(n2746), .B(n1710), .Z(o_m_imm[0]) );
  HDOAI211D1 U2317 ( .A1(n2956), .A2(n1732), .B(n2955), .C(n2954), .Z(n2957)
         );
  HDOAI22D1 U2318 ( .A1(n2948), .A2(n2814), .B1(n2813), .B2(n2810), .Z(
        o_rs1[2]) );
  HDOAI211D1 U2319 ( .A1(n2805), .A2(n2939), .B(n2804), .C(n2803), .Z(n2806)
         );
  HDINVD1 U2320 ( .A(n2802), .Z(n2803) );
  HDAOI21D1 U2321 ( .A1(n2881), .A2(n1767), .B(n1766), .Z(n2961) );
  HDNAN4D1 U2322 ( .A1(n2707), .A2(n412), .A3(n410), .A4(n1765), .Z(n1767) );
  HDNAN2D1 U2323 ( .A1(n1764), .A2(n2899), .Z(n1765) );
  HDOAI211D1 U2324 ( .A1(n1897), .A2(n1902), .B(n1709), .C(n1896), .Z(
        o_m_imm[4]) );
  HDNAN2D1 U2325 ( .A1(n1926), .A2(o_rs2_2_), .Z(n1896) );
  HDNAN2D1 U2326 ( .A1(n2833), .A2(n2832), .Z(o_rd2[0]) );
  HDOAI211D1 U2327 ( .A1(n1897), .A2(n1998), .B(n1905), .C(n1895), .Z(
        o_m_imm[3]) );
  HDNAN2D1 U2328 ( .A1(n1926), .A2(o_rs2_1_), .Z(n1895) );
  HDOAI211D1 U2329 ( .A1(n1907), .A2(n2979), .B(n1904), .C(n1710), .Z(
        o_m_imm[8]) );
  HDNAN2D1 U2330 ( .A1(n1926), .A2(instruction[6]), .Z(n1904) );
  HDOAI211D1 U2331 ( .A1(n1907), .A2(n2980), .B(n1903), .C(n1709), .Z(
        o_m_imm[7]) );
  HDNAN2D1 U2332 ( .A1(n1926), .A2(instruction[5]), .Z(n1903) );
  HDOAI211D1 U2333 ( .A1(n1907), .A2(n1947), .B(n1906), .C(n1905), .Z(
        o_m_imm[9]) );
  HDNAN2D1 U2334 ( .A1(n1926), .A2(instruction[7]), .Z(n1906) );
  HDOAI21D1 U2335 ( .A1(n2638), .A2(n1732), .B(n2637), .Z(o_rs4[5]) );
  HDNOR4D1 U2336 ( .A1(n2848), .A2(n2636), .A3(n2635), .A4(n2634), .Z(n2638)
         );
  HDAOI31D1 U2337 ( .A1(n2631), .A2(n2630), .A3(n2629), .B(n2628), .Z(n2636)
         );
  HDINVD1 U2338 ( .A(n2622), .Z(n2623) );
  HDINVD1 U2339 ( .A(n1717), .Z(n1718) );
  HDAOI21D1 U2340 ( .A1(n1732), .A2(n2489), .B(n2488), .Z(o_m_futype[1]) );
  HDNOR4D1 U2341 ( .A1(n2487), .A2(n2486), .A3(n2485), .A4(n2484), .Z(n2488)
         );
  HDOAI22D1 U2342 ( .A1(n2929), .A2(n2927), .B1(n2480), .B2(n835), .Z(n2485)
         );
  HDINVD1 U2343 ( .A(n2967), .Z(n2480) );
  HDOAI31D1 U2344 ( .A1(n2523), .A2(n2522), .A3(n2478), .B(n1599), .Z(n2489)
         );
  HDAND2D1 U2345 ( .A1(n2824), .A2(n1744), .Z(n2832) );
  HDINVD1 U2346 ( .A(o_m_flags[3]), .Z(n1744) );
  HDNOR2D1 U2347 ( .A1(n2815), .A2(n1732), .Z(o_rd2_type[3]) );
  HDINVD1 U2348 ( .A(n2333), .Z(n2815) );
  HDAOI22D1 U2349 ( .A1(instruction[16]), .A2(n2687), .B1(n2686), .B2(n2685), 
        .Z(n2689) );
  HDAO211D1 U2350 ( .A1(n2230), .A2(n1609), .B(n2497), .C(n2229), .Z(
        o_m_opcode[2]) );
  HDOAI22D1 U2351 ( .A1(n2228), .A2(n1737), .B1(n2227), .B2(n2934), .Z(n2229)
         );
  HDNOR4D1 U2352 ( .A1(n2226), .A2(n2225), .A3(n2224), .A4(n2223), .Z(n2227)
         );
  HDNAN3D1 U2353 ( .A1(n2432), .A2(n2208), .A3(n2207), .Z(n2226) );
  HDNOR4D1 U2354 ( .A1(n2206), .A2(n2205), .A3(n2204), .A4(n2203), .Z(n2228)
         );
  HDINVD1 U2355 ( .A(n2200), .Z(n2201) );
  HDNAN4D1 U2356 ( .A1(n2197), .A2(n2196), .A3(n2195), .A4(n2194), .Z(n2230)
         );
  HDNOR4D1 U2357 ( .A1(n2193), .A2(n2192), .A3(n2406), .A4(n2585), .Z(n2194)
         );
  HDNAN3D1 U2358 ( .A1(n2268), .A2(n2251), .A3(n2328), .Z(n2193) );
  HDAOI211D1 U2359 ( .A1(n2685), .A2(n2795), .B(n2429), .C(n2181), .Z(n2195)
         );
  HDOAI211D1 U2360 ( .A1(n2180), .A2(n2443), .B(n2179), .C(n2178), .Z(n2181)
         );
  HDAOI211D1 U2361 ( .A1(n2360), .A2(n2173), .B(n2172), .C(n2645), .Z(n2196)
         );
  HDAOI211D1 U2362 ( .A1(n2169), .A2(n2881), .B(n2168), .C(n2167), .Z(n2197)
         );
  HDAOI21D1 U2363 ( .A1(n1619), .A2(n2160), .B(n2417), .Z(n2168) );
  HDAND2D1 U2364 ( .A1(n2975), .A2(n2899), .Z(n472) );
  HDOAI211D1 U2365 ( .A1(n2595), .A2(n1737), .B(n2637), .C(n2594), .Z(o_rs4[2]) );
  HDOAI31D1 U2366 ( .A1(n2593), .A2(n2839), .A3(n2634), .B(n1609), .Z(n2594)
         );
  HDOAI22D1 U2367 ( .A1(n2588), .A2(n2628), .B1(n2603), .B2(n2614), .Z(n2593)
         );
  HDNOR2D1 U2368 ( .A1(n2556), .A2(n2555), .Z(n2557) );
  HDINVD1 U2369 ( .A(n2614), .Z(n2555) );
  HDNOR4D1 U2370 ( .A1(n2587), .A2(n2586), .A3(n2585), .A4(n2584), .Z(n2595)
         );
  HDNAN4D1 U2371 ( .A1(n2583), .A2(n2873), .A3(n2582), .A4(n2581), .Z(n2584)
         );
  HDOAI222D1 U2372 ( .A1(n1737), .A2(n2433), .B1(n2934), .B2(n2432), .C1(n1732), .C2(n2431), .Z(o_m_opcode[7]) );
  HDNOR4D1 U2373 ( .A1(n2430), .A2(n2429), .A3(n2428), .A4(n2427), .Z(n2431)
         );
  HDOAI21D1 U2374 ( .A1(n2426), .A2(n2425), .B(n2424), .Z(n2427) );
  HDOAI211D1 U2375 ( .A1(n2423), .A2(n2422), .B(n2421), .C(n2420), .Z(n2428)
         );
  HDINVD1 U2376 ( .A(n2445), .Z(n2420) );
  HDNAN4D1 U2377 ( .A1(n2419), .A2(n2418), .A3(n2417), .A4(n2416), .Z(n2430)
         );
  HDNOR3D1 U2378 ( .A1(n2414), .A2(n2413), .A3(n2412), .Z(n2419) );
  HDINVD1 U2379 ( .A(n2411), .Z(n2413) );
  HDAOI21D1 U2380 ( .A1(n2241), .A2(n2373), .B(n2257), .Z(n2432) );
  HDINVD1 U2381 ( .A(n2521), .Z(n2410) );
  HDNAN2D1 U2382 ( .A1(n1612), .A2(n2457), .Z(o_m_opcode[8]) );
  HDNOR2D1 U2383 ( .A1(n2440), .A2(n1614), .Z(n2449) );
  HDOR3D1 U2384 ( .A1(n2750), .A2(n2438), .A3(n2439), .Z(n1614) );
  HDINVD1 U2385 ( .A(n2434), .Z(n2440) );
  HDOAI21D1 U2386 ( .A1(n2455), .A2(n2454), .B(n1599), .Z(n2456) );
  HDOAI211D1 U2387 ( .A1(n1828), .A2(n1732), .B(n1827), .C(n1826), .Z(o_fail)
         );
  HDNOR3D1 U2388 ( .A1(n1704), .A2(n2678), .A3(n2934), .Z(n1871) );
  HDNOR4D1 U2389 ( .A1(n1818), .A2(n1817), .A3(n1816), .A4(n1815), .Z(n1828)
         );
  HDOAI222D1 U2390 ( .A1(n2930), .A2(n1814), .B1(n2359), .B2(n1806), .C1(n2679), .C2(n1813), .Z(n1815) );
  HDNOR3D1 U2391 ( .A1(n1810), .A2(n1702), .A3(n1809), .Z(n1814) );
  HDOAI211D1 U2392 ( .A1(n2063), .A2(n2062), .B(n1808), .C(n2742), .Z(n1810)
         );
  HDINVD1 U2393 ( .A(n2923), .Z(n1808) );
  HDNOR2D1 U2394 ( .A1(n2447), .A2(n2356), .Z(n1875) );
  HDAOI211D1 U2395 ( .A1(n2976), .A2(n1799), .B(n1550), .C(n1798), .Z(n1805)
         );
  HDINVD1 U2396 ( .A(n2718), .Z(n1799) );
  HDOAI211D1 U2397 ( .A1(n1623), .A2(n1732), .B(n1624), .C(n1600), .Z(
        o_m_opcode[4]) );
  HDAOI22D1 U2398 ( .A1(n2941), .A2(n1625), .B1(n1626), .B2(n1599), .Z(n1624)
         );
  HDINVD1 U2399 ( .A(n2328), .Z(n1627) );
  HDNOR2D1 U2400 ( .A1(n2384), .A2(n2191), .Z(n2328) );
  HDNOR2D1 U2401 ( .A1(n1632), .A2(n1610), .Z(n1623) );
  HDOR2D1 U2402 ( .A1(n1634), .A2(n1633), .Z(n1610) );
  HDOAI211D1 U2403 ( .A1(instruction[5]), .A2(n2320), .B(n2421), .C(n1635), 
        .Z(n1633) );
  HDAOI21D1 U2404 ( .A1(n2387), .A2(n2443), .B(n2389), .Z(n1636) );
  HDNAN4D1 U2405 ( .A1(n2434), .A2(n1637), .A3(n2344), .A4(n2390), .Z(n1632)
         );
  HDAND4D1 U2406 ( .A1(n2306), .A2(n2385), .A3(n1621), .A4(n2307), .Z(n2434)
         );
  HDINVD1 U2407 ( .A(n2308), .Z(n2426) );
  HDOAI211D1 U2408 ( .A1(n1936), .A2(n2977), .B(n1935), .C(n1938), .Z(
        o_m_imm[15]) );
  HDNAN2D1 U2409 ( .A1(n2876), .A2(instruction[5]), .Z(n1935) );
  HDOAI211D1 U2410 ( .A1(n1936), .A2(n2064), .B(n1933), .C(n1938), .Z(
        o_m_imm[13]) );
  HDNAN2D1 U2411 ( .A1(n2876), .A2(o_rs2_3_), .Z(n1933) );
  HDOAI211D1 U2412 ( .A1(n1932), .A2(n1931), .B(n1930), .C(n1938), .Z(
        o_m_imm[12]) );
  HDAOI22D1 U2413 ( .A1(n2876), .A2(o_rs2_2_), .B1(n1926), .B2(instruction[10]), .Z(n1930) );
  HDINVD1 U2414 ( .A(n1927), .Z(n1931) );
  HDINVD1 U2415 ( .A(n2506), .Z(n1932) );
  HDOAI211D1 U2416 ( .A1(n1936), .A2(n2399), .B(n1934), .C(n1938), .Z(
        o_m_imm[14]) );
  HDNAN2D1 U2417 ( .A1(n2876), .A2(o_rs2_4_), .Z(n1934) );
  HDOAI211D1 U2418 ( .A1(n1940), .A2(n2797), .B(n1939), .C(n1938), .Z(
        o_m_imm[16]) );
  HDAOI22D1 U2419 ( .A1(instruction[20]), .A2(n2770), .B1(n2876), .B2(
        instruction[6]), .Z(n1939) );
  HDINVD1 U2420 ( .A(n1948), .Z(n1940) );
  HDOAI21D1 U2421 ( .A1(n2592), .A2(n2604), .B(n2591), .Z(n2839) );
  HDNOR2D1 U2422 ( .A1(n1793), .A2(n2929), .Z(n424) );
  HDAOI211D1 U2423 ( .A1(n1792), .A2(n2899), .B(n2896), .C(n1791), .Z(n1793)
         );
  HDOAI211D1 U2424 ( .A1(n2709), .A2(n2902), .B(n412), .C(n1790), .Z(n1791) );
  HDINVD1 U2425 ( .A(n457), .Z(n1792) );
  HDOAI211D1 U2426 ( .A1(n2519), .A2(n1737), .B(n2518), .C(n2517), .Z(
        o_m_type[0]) );
  HDNAN2D1 U2427 ( .A1(n2516), .A2(n1735), .Z(n2517) );
  HDOAI211D1 U2428 ( .A1(n2515), .A2(n2604), .B(n2514), .C(n2513), .Z(n2516)
         );
  HDNOR3D1 U2429 ( .A1(n2512), .A2(n2883), .A3(n1652), .Z(n2513) );
  HDAOI22D1 U2430 ( .A1(n2941), .A2(n2453), .B1(n2452), .B2(n1599), .Z(n2518)
         );
  HDNOR4D1 U2431 ( .A1(n2523), .A2(n2778), .A3(n2499), .A4(n2498), .Z(n2519)
         );
  HDINVD1 U2432 ( .A(n2733), .Z(n2498) );
  HDOAI211D1 U2433 ( .A1(n2613), .A2(n1732), .B(n2637), .C(n2836), .Z(o_rs4[3]) );
  HDNOR4D1 U2434 ( .A1(n2612), .A2(n2611), .A3(n2842), .A4(n2610), .Z(n2613)
         );
  HDOAI211D1 U2435 ( .A1(n2952), .A2(n2819), .B(n2609), .C(n2608), .Z(n2842)
         );
  HDAOI211D1 U2436 ( .A1(n2607), .A2(n2981), .B(n2622), .C(n2606), .Z(n2608)
         );
  HDNOR2D1 U2437 ( .A1(n2605), .A2(n2604), .Z(n2606) );
  HDOAI211D1 U2438 ( .A1(n2603), .A2(n2602), .B(n2601), .C(n2600), .Z(n2612)
         );
  HDINVD1 U2439 ( .A(n2559), .Z(n2596) );
  HDOAI211D1 U2440 ( .A1(n1936), .A2(n1902), .B(n1905), .C(n1901), .Z(
        o_m_imm[6]) );
  HDNAN2D1 U2441 ( .A1(n1900), .A2(instruction[6]), .Z(n1901) );
  HDINVD1 U2442 ( .A(o_rs2_4_), .Z(n1902) );
  HDOAI211D1 U2443 ( .A1(n1859), .A2(n1737), .B(n1858), .C(n1857), .Z(
        o_m_flags[6]) );
  HDNOR4D1 U2444 ( .A1(n2547), .A2(n2845), .A3(n2834), .A4(n2590), .Z(n1854)
         );
  HDNOR3D1 U2445 ( .A1(n2849), .A2(n1837), .A3(n2533), .Z(n1858) );
  HDNOR3D1 U2446 ( .A1(n1836), .A2(n2406), .A3(n2407), .Z(n1859) );
  HDAOI22D1 U2447 ( .A1(n2795), .A2(instruction[25]), .B1(n2794), .B2(
        instruction[14]), .Z(n2796) );
  HDOAI211D1 U2448 ( .A1(n2793), .A2(n2929), .B(n2792), .C(n2791), .Z(n2794)
         );
  HDNOR2D1 U2449 ( .A1(n2808), .A2(n2790), .Z(n2791) );
  HDNOR4D1 U2450 ( .A1(n2788), .A2(n2787), .A3(n2878), .A4(n2786), .Z(n2793)
         );
  HDNOR3D1 U2451 ( .A1(n2852), .A2(n2976), .A3(n2979), .Z(n919) );
  HDNOR2D1 U2452 ( .A1(n2953), .A2(n2952), .Z(o_rd[4]) );
  HDNAN2D1 U2453 ( .A1(n1618), .A2(n2888), .Z(n2890) );
  HDAOI22M10D1 U2454 ( .B1(n2894), .B2(n2911), .A1(n1724), .A2(n2881), .Z(
        n2888) );
  HDOA21M20D1 U2455 ( .A1(n2878), .A2(n2974), .B(n631), .Z(n1724) );
  HDNAN2D1 U2456 ( .A1(n2927), .A2(n2415), .Z(n2878) );
  HDAOI211D1 U2457 ( .A1(n2886), .A2(n2973), .B(n2885), .C(n2884), .Z(n2887)
         );
  HDNAN2D1 U2458 ( .A1(n2355), .A2(n395), .Z(n2882) );
  HDNAN2D1 U2459 ( .A1(n2852), .A2(n2901), .Z(n2886) );
  HDOAI211D1 U2460 ( .A1(n2693), .A2(n2809), .B(n2684), .C(n2683), .Z(o_rs3[1]) );
  HDAOI21D1 U2461 ( .A1(n2691), .A2(instruction[26]), .B(n2682), .Z(n2683) );
  HDINVD1 U2462 ( .A(instruction[20]), .Z(n2678) );
  HDOAI211D1 U2463 ( .A1(instruction[11]), .A2(instruction[12]), .B(n2675), 
        .C(n2686), .Z(n2684) );
  HDINVD1 U2464 ( .A(n360), .Z(n2686) );
  HDNAN2D1 U2465 ( .A1(n2909), .A2(n1735), .Z(n2910) );
  HDAOI211D1 U2466 ( .A1(n2906), .A2(n2905), .B(n2904), .C(n2903), .Z(n2956)
         );
  HDOAI22D1 U2467 ( .A1(n2902), .A2(n2901), .B1(n2900), .B2(n2929), .Z(n2904)
         );
  HDAOI211D1 U2468 ( .A1(n2899), .A2(n590), .B(n2898), .C(n2897), .Z(n2900) );
  HDNAN2M1D1 U2469 ( .A1(n2896), .A2(n2895), .Z(n2898) );
  HDNOR2M1D1 U2470 ( .A1(n599), .A2(n2987), .Z(n2896) );
  HDNAN2D1 U2471 ( .A1(n388), .A2(n457), .Z(n599) );
  HDNAN2D1 U2472 ( .A1(n2725), .A2(n2979), .Z(n457) );
  HDNAN2M1D1 U2473 ( .A1(n2880), .A2(n2879), .Z(n2894) );
  HDNOR4D1 U2474 ( .A1(n2861), .A2(n2860), .A3(n2859), .A4(n2858), .Z(n2879)
         );
  HDNAN2D1 U2475 ( .A1(n2892), .A2(n1599), .Z(n2955) );
  HDAOI21D1 U2476 ( .A1(n2877), .A2(n1599), .B(n2876), .Z(n2912) );
  HDOAI211D1 U2477 ( .A1(n2746), .A2(n2868), .B(n1918), .C(n1917), .Z(
        o_m_imm[10]) );
  HDAOI211D1 U2478 ( .A1(instruction[8]), .A2(n1926), .B(n1728), .C(n1916), 
        .Z(n1917) );
  HDNOR4D1 U2479 ( .A1(n2367), .A2(n2366), .A3(n2365), .A4(n2364), .Z(n2368)
         );
  HDOAI211D1 U2480 ( .A1(n2363), .A2(n2976), .B(n2362), .C(n2361), .Z(n2364)
         );
  HDNOR2D1 U2481 ( .A1(n2866), .A2(n2644), .Z(n2362) );
  HDOAI211D1 U2482 ( .A1(n2394), .A2(n2359), .B(n2358), .C(n2357), .Z(n2365)
         );
  HDNAN3D1 U2483 ( .A1(n2351), .A2(n2350), .A3(n2349), .Z(n2366) );
  HDINVD1 U2484 ( .A(n2346), .Z(n2347) );
  HDINVD1 U2485 ( .A(n2469), .Z(n2351) );
  HDNOR2D1 U2486 ( .A1(n399), .A2(n2980), .Z(n2469) );
  HDNAN3D1 U2487 ( .A1(n2345), .A2(n2344), .A3(n2343), .Z(n2367) );
  HDAOI211D1 U2488 ( .A1(n922), .A2(n2723), .B(n593), .C(n2314), .Z(n2316) );
  HDNOR3D1 U2489 ( .A1(n2342), .A2(n2341), .A3(n2412), .Z(n2345) );
  HDNAN4D1 U2490 ( .A1(n2442), .A2(n2436), .A3(n2390), .A4(n2386), .Z(n2412)
         );
  HDINVD1 U2491 ( .A(n2483), .Z(n2341) );
  HDNOR4D1 U2492 ( .A1(n2371), .A2(n2335), .A3(n2334), .A4(n2333), .Z(n2370)
         );
  HDNAN2D1 U2493 ( .A1(n2872), .A2(n2673), .Z(n2333) );
  HDNAN3D1 U2494 ( .A1(n2332), .A2(n2738), .A3(n2604), .Z(n2334) );
  HDOAI22D1 U2495 ( .A1(n2812), .A2(n2693), .B1(n2692), .B2(n2952), .Z(
        o_rs3[4]) );
  HDOAI22D1 U2496 ( .A1(n2811), .A2(n2693), .B1(n2692), .B2(n2951), .Z(
        o_rs3[3]) );
  HDINVD1 U2497 ( .A(n2691), .Z(n2692) );
  HDAOI21D1 U2498 ( .A1(n2677), .A2(n2676), .B(n1736), .Z(n2691) );
  HDOAI211D1 U2499 ( .A1(n2754), .A2(n1732), .B(n2753), .C(n475), .Z(
        o_rs1_valid) );
  HDNAN2D1 U2500 ( .A1(n1757), .A2(n1599), .Z(n475) );
  HDNOR3D1 U2501 ( .A1(n2455), .A2(n2522), .A3(n2920), .Z(n1755) );
  HDNAN4D1 U2502 ( .A1(n1754), .A2(n2044), .A3(n2493), .A4(n2267), .Z(n2455)
         );
  HDINVD1 U2503 ( .A(n1863), .Z(n1756) );
  HDAND4D1 U2504 ( .A1(n2752), .A2(n2751), .A3(n2962), .A4(n2798), .Z(n2754)
         );
  HDNOR2D1 U2505 ( .A1(n1766), .A2(n488), .Z(n2962) );
  HDAOI21D1 U2506 ( .A1(n1762), .A2(n2852), .B(n2853), .Z(n1766) );
  HDNOR4D1 U2507 ( .A1(n2750), .A2(n2749), .A3(n2862), .A4(n2748), .Z(n2752)
         );
  HDNAN3D1 U2508 ( .A1(n2530), .A2(n2436), .A3(n2767), .Z(n2750) );
  HDINVD1 U2509 ( .A(n2773), .Z(n2436) );
  HDNAN2D1 U2510 ( .A1(n2824), .A2(n2553), .Z(o_rs4[0]) );
  HDOAI31D1 U2511 ( .A1(n2552), .A2(n2610), .A3(n2831), .B(n1609), .Z(n2553)
         );
  HDOAI211D1 U2512 ( .A1(n2551), .A2(n2550), .B(n2569), .C(n2549), .Z(n2831)
         );
  HDNOR2D1 U2513 ( .A1(n2622), .A2(n2547), .Z(n2569) );
  HDNOR2D1 U2514 ( .A1(n2546), .A2(n2551), .Z(n2622) );
  HDOAI22M10D1 U2515 ( .A1(n2545), .A2(n2603), .B1(n2544), .B2(n2628), .Z(
        n2552) );
  HDNOR4D1 U2516 ( .A1(n2554), .A2(n2561), .A3(n2540), .A4(n2539), .Z(n2598)
         );
  HDNAN3D1 U2517 ( .A1(n2537), .A2(instruction[14]), .A3(n2536), .Z(n2614) );
  HDINVD1 U2518 ( .A(n2535), .Z(n2616) );
  HDAND2D1 U2519 ( .A1(n2840), .A2(n2836), .Z(n2824) );
  HDOAI211D1 U2520 ( .A1(n2580), .A2(n2977), .B(n2375), .C(n1742), .Z(n2836)
         );
  HDNOR2D1 U2521 ( .A1(n2987), .A2(n1442), .Z(n2580) );
  HDNAN4D1 U2522 ( .A1(o_rs2_2_), .A2(n2971), .A3(o_rs2_4_), .A4(n1443), .Z(
        n1442) );
  HDNAN2D1 U2523 ( .A1(n1789), .A2(n1788), .Z(n528) );
  HDOAI22D1 U2524 ( .A1(n388), .A2(n2696), .B1(n1786), .B2(n2797), .Z(n1789)
         );
  HDNOR2D1 U2525 ( .A1(n1787), .A2(n2725), .Z(n1786) );
  HDOAI211D1 U2526 ( .A1(n2916), .A2(n2744), .B(n2775), .C(n1785), .Z(n1787)
         );
  HDINVD1 U2527 ( .A(n2903), .Z(n1785) );
  HDNAN3D1 U2528 ( .A1(n2963), .A2(n2774), .A3(n2387), .Z(n2903) );
  HDNOR2D1 U2529 ( .A1(n2611), .A2(n2773), .Z(n2963) );
  HDOAI211D1 U2530 ( .A1(n1936), .A2(n1998), .B(n1709), .C(n1899), .Z(
        o_m_imm[5]) );
  HDOAI21D1 U2531 ( .A1(n1900), .A2(n1927), .B(instruction[5]), .Z(n1899) );
  HDOAI22D1 U2532 ( .A1(n2772), .A2(n1732), .B1(n2782), .B2(n2771), .Z(
        o_rs1_type[0]) );
  HDNOR3D1 U2533 ( .A1(n2758), .A2(n2757), .A3(n2756), .Z(n2772) );
  HDINVD1 U2534 ( .A(n1615), .Z(o_m_imm_44_) );
  HDINVD1 U2535 ( .A(n1615), .Z(o_m_imm_40_) );
  HDINVD1 U2536 ( .A(n1615), .Z(o_m_imm_38_) );
  HDINVD1 U2537 ( .A(n1615), .Z(o_m_imm_52_) );
  HDAOI22D1 U2538 ( .A1(instruction[22]), .A2(n2497), .B1(n2876), .B2(
        instruction[14]), .Z(n1957) );
  HDAOI22D1 U2539 ( .A1(n2497), .A2(instruction[26]), .B1(n2876), .B2(
        instruction[18]), .Z(n1961) );
  HDAOI22D1 U2540 ( .A1(n2497), .A2(instruction[27]), .B1(n2876), .B2(
        instruction[19]), .Z(n1962) );
  HDAOI22D1 U2541 ( .A1(instruction[21]), .A2(n2497), .B1(n2876), .B2(
        instruction[13]), .Z(n1956) );
  HDAOI22D1 U2542 ( .A1(instruction[23]), .A2(n2497), .B1(n2876), .B2(
        instruction[15]), .Z(n1958) );
  HDAOI22D1 U2543 ( .A1(instruction[25]), .A2(n2497), .B1(n2876), .B2(
        instruction[17]), .Z(n1960) );
  HDAOI22D1 U2544 ( .A1(instruction[24]), .A2(n2497), .B1(n2876), .B2(
        instruction[16]), .Z(n1959) );
  HDAOI22D1 U2545 ( .A1(n2497), .A2(instruction[28]), .B1(n2876), .B2(
        instruction[20]), .Z(n1963) );
  HDNAN2D1 U2546 ( .A1(n1703), .A2(n2302), .Z(o_m_opcode[3]) );
  HDNAN4D1 U2547 ( .A1(n2300), .A2(n2299), .A3(n2298), .A4(n2297), .Z(n2301)
         );
  HDNOR2D1 U2548 ( .A1(n2901), .A2(n2290), .Z(n2293) );
  HDINVD1 U2549 ( .A(n2713), .Z(n2290) );
  HDNAN2D1 U2550 ( .A1(n2163), .A2(n2675), .Z(n2294) );
  HDOR2D1 U2551 ( .A1(instruction[15]), .A2(instruction[16]), .Z(n1619) );
  HDINVD1 U2552 ( .A(n2318), .Z(n2447) );
  HDAOI211D1 U2553 ( .A1(n990), .A2(n2481), .B(n2280), .C(n2279), .Z(n2299) );
  HDOAI22D1 U2554 ( .A1(n2278), .A2(n2767), .B1(n2852), .B2(n2277), .Z(n2279)
         );
  HDNOR2D1 U2555 ( .A1(n2273), .A2(n1613), .Z(n2300) );
  HDOR3D1 U2556 ( .A1(n2272), .A2(n2340), .A3(n2441), .Z(n1613) );
  HDAND2D1 U2557 ( .A1(n2966), .A2(n2881), .Z(n488) );
  HDINVD1 U2558 ( .A(n2834), .Z(n2267) );
  HDAOI211D1 U2559 ( .A1(n2188), .A2(n2883), .B(n2315), .C(n2187), .Z(n2268)
         );
  HDNAN2D1 U2560 ( .A1(n2185), .A2(n2184), .Z(n2188) );
  HDNOR2D1 U2561 ( .A1(n2414), .A2(n2572), .Z(n2269) );
  HDINVD1 U2562 ( .A(n2530), .Z(n2414) );
  HDNOR2D1 U2563 ( .A1(n2263), .A2(n2527), .Z(n2411) );
  HDOA21D1 U2564 ( .A1(n2304), .A2(n2934), .B(n2303), .Z(n1703) );
  HDOAI21D1 U2565 ( .A1(n2262), .A2(n2261), .B(n1599), .Z(n2303) );
  HDINVD1 U2566 ( .A(n2454), .Z(n2253) );
  HDOR2D1 U2567 ( .A1(n2733), .A2(instruction[0]), .Z(n2332) );
  HDINVD1 U2568 ( .A(n2478), .Z(n2873) );
  HDNOR3D1 U2569 ( .A1(n2329), .A2(n2870), .A3(n2252), .Z(n2255) );
  HDNOR4D1 U2570 ( .A1(n2190), .A2(n2522), .A3(n2441), .A4(n2200), .Z(n2251)
         );
  HDNAN2D1 U2571 ( .A1(n2331), .A2(n2349), .Z(n2190) );
  HDNOR4D1 U2572 ( .A1(n2250), .A2(n2249), .A3(n2248), .A4(n2247), .Z(n2304)
         );
  HDOAI211D1 U2573 ( .A1(n2278), .A2(n1704), .B(n2239), .C(n2238), .Z(n2250)
         );
  HDOAI21D1 U2574 ( .A1(n2237), .A2(n2236), .B(n2235), .Z(n2238) );
  HDNAN2D1 U2575 ( .A1(n2215), .A2(n2209), .Z(n2237) );
  HDNOR2D1 U2576 ( .A1(n2232), .A2(n2339), .Z(n2278) );
  HDNAN3D1 U2577 ( .A1(n2802), .A2(n1735), .A3(instruction[14]), .Z(n2695) );
  HDAOI21D1 U2578 ( .A1(n2653), .A2(n2798), .B(n1732), .Z(n2687) );
  HDINVD1 U2579 ( .A(o_rd_type[3]), .Z(n2954) );
  HDOAI211D1 U2580 ( .A1(n2672), .A2(n1732), .B(n2671), .C(n2670), .Z(
        o_rs3_type[1]) );
  HDNOR4D1 U2581 ( .A1(n2645), .A2(n2644), .A3(n2643), .A4(n2642), .Z(n2647)
         );
  HDNOR2D1 U2582 ( .A1(n2854), .A2(n2976), .Z(n2643) );
  HDNAN2D1 U2583 ( .A1(n2639), .A2(n2980), .Z(n2854) );
  HDNAN2D1 U2584 ( .A1(n2669), .A2(n1599), .Z(n2671) );
  HDINVD1 U2585 ( .A(n2920), .Z(n2657) );
  HDAOI21D1 U2586 ( .A1(n2665), .A2(n2771), .B(n2664), .Z(n2672) );
  HDNOR2D1 U2587 ( .A1(n2099), .A2(n2795), .Z(n2663) );
  HDINVD1 U2588 ( .A(n1615), .Z(o_m_imm_48_) );
  HDINVD1 U2589 ( .A(n1615), .Z(o_m_imm_42_) );
  HDNOR3D1 U2590 ( .A1(n1971), .A2(n1970), .A3(n1969), .Z(n1972) );
  HDINVD1 U2591 ( .A(n1728), .Z(n1973) );
  HDOAI211D1 U2592 ( .A1(n2405), .A2(n2934), .B(n2404), .C(n2403), .Z(
        o_m_opcode[6]) );
  HDOAI31D1 U2593 ( .A1(n2402), .A2(n2401), .A3(n2400), .B(n1609), .Z(n2403)
         );
  HDOAI211D1 U2594 ( .A1(n2918), .A2(n2399), .B(n2398), .C(n2397), .Z(n2400)
         );
  HDNOR2D1 U2595 ( .A1(n2929), .A2(n2976), .Z(n2967) );
  HDOAI211D1 U2596 ( .A1(n2396), .A2(n2929), .B(n2395), .C(n2424), .Z(n2401)
         );
  HDOR2D1 U2597 ( .A1(n2653), .A2(n2394), .Z(n2424) );
  HDNOR2D1 U2598 ( .A1(instruction[10]), .A2(instruction[11]), .Z(n2394) );
  HDNAN3D1 U2599 ( .A1(n2800), .A2(instruction[7]), .A3(n387), .Z(n2653) );
  HDINVD1 U2600 ( .A(n2390), .Z(n2391) );
  HDOR2D1 U2601 ( .A1(n2318), .A2(n2446), .Z(n2390) );
  HDOR2D1 U2602 ( .A1(n2317), .A2(instruction[16]), .Z(n2446) );
  HDNAN2D1 U2603 ( .A1(n2505), .A2(instruction[18]), .Z(n2318) );
  HDINVD1 U2604 ( .A(n2352), .Z(n2389) );
  HDNOR2D1 U2605 ( .A1(n2310), .A2(n2811), .Z(n2352) );
  HDINVD1 U2606 ( .A(n2639), .Z(n2393) );
  HDAND2D1 U2607 ( .A1(n2313), .A2(n2312), .Z(n2396) );
  HDNAN2D1 U2608 ( .A1(n2158), .A2(n1094), .Z(n2312) );
  HDAOI21D1 U2609 ( .A1(n2899), .A2(n2291), .B(n2964), .Z(n2313) );
  HDNAN2D1 U2610 ( .A1(n647), .A2(n671), .Z(n2291) );
  HDNAN4D1 U2611 ( .A1(n2388), .A2(n2632), .A3(n2387), .A4(n2386), .Z(n2402)
         );
  HDINVD1 U2612 ( .A(n2340), .Z(n2386) );
  HDAOI21D1 U2613 ( .A1(n2270), .A2(n2538), .B(n2443), .Z(n2340) );
  HDNAN2D1 U2614 ( .A1(n2639), .A2(n2799), .Z(n2387) );
  HDAOI222D1 U2615 ( .A1(n2381), .A2(n1599), .B1(n2380), .B2(n2646), .C1(n2379), .C2(n2378), .Z(n2404) );
  HDNOR2D1 U2616 ( .A1(n2753), .A2(instruction[28]), .Z(n2378) );
  HDINVD1 U2617 ( .A(n2493), .Z(n2666) );
  HDOAI211D1 U2618 ( .A1(n1936), .A2(n2746), .B(n1710), .C(n1894), .Z(
        o_m_imm[2]) );
  HDNAN2D1 U2619 ( .A1(n1893), .A2(o_rs2_2_), .Z(n1894) );
  HDNOR3D1 U2620 ( .A1(n1912), .A2(n2883), .A3(n1910), .Z(n1887) );
  HDOAI211D1 U2621 ( .A1(n2868), .A2(n2979), .B(n1945), .C(n1949), .Z(
        o_m_imm[18]) );
  HDNAN2D1 U2622 ( .A1(n1948), .A2(instruction[16]), .Z(n1945) );
  HDOAI211D1 U2623 ( .A1(n2868), .A2(n2980), .B(n1944), .C(n1949), .Z(
        o_m_imm[17]) );
  HDNAN2D1 U2624 ( .A1(n1948), .A2(instruction[15]), .Z(n1944) );
  HDOAI211D1 U2625 ( .A1(n2868), .A2(n1947), .B(n1946), .C(n1949), .Z(
        o_m_imm[19]) );
  HDNAN2D1 U2626 ( .A1(n1948), .A2(instruction[17]), .Z(n1946) );
  HDOAI211D1 U2627 ( .A1(n2868), .A2(n2978), .B(n1950), .C(n1949), .Z(
        o_m_imm[20]) );
  HDINVD1 U2628 ( .A(n1953), .Z(n1943) );
  HDNAN2D1 U2629 ( .A1(n1948), .A2(instruction[18]), .Z(n1950) );
  HDNAN2D1 U2630 ( .A1(n1937), .A2(n1600), .Z(n1948) );
  HDOAI211D1 U2631 ( .A1(n2157), .A2(n1732), .B(n2156), .C(n1600), .Z(
        o_m_opcode[1]) );
  HDAOI22M10D1 U2632 ( .B1(n2155), .B2(n1599), .A1(n2154), .A2(n2941), .Z(
        n2156) );
  HDNAN4D1 U2633 ( .A1(n2208), .A2(n2151), .A3(n2150), .A4(n2149), .Z(n2152)
         );
  HDNOR2D1 U2634 ( .A1(n2379), .A2(n2948), .Z(n2211) );
  HDINVD1 U2635 ( .A(n2453), .Z(n2151) );
  HDNAN2D1 U2636 ( .A1(n2215), .A2(n2321), .Z(n2144) );
  HDNAN2D1 U2637 ( .A1(n2339), .A2(n2951), .Z(n2215) );
  HDNAN4D1 U2638 ( .A1(n2143), .A2(n2142), .A3(n2654), .A4(n2331), .Z(n2155)
         );
  HDNAN2D1 U2639 ( .A1(n2179), .A2(n2140), .Z(n2141) );
  HDNAN2D1 U2640 ( .A1(n2139), .A2(n2501), .Z(n2179) );
  HDNAN2D1 U2641 ( .A1(n1687), .A2(n2199), .Z(n2139) );
  HDNOR2D1 U2642 ( .A1(n1720), .A2(n2659), .Z(n2667) );
  HDNOR3D1 U2643 ( .A1(n2138), .A2(n2137), .A3(n2136), .Z(n2143) );
  HDINVD1 U2644 ( .A(n2451), .Z(n2137) );
  HDNOR2D1 U2645 ( .A1(n2749), .A2(n2200), .Z(n2451) );
  HDNOR4D1 U2646 ( .A1(n2135), .A2(n2134), .A3(n2133), .A4(n2132), .Z(n2157)
         );
  HDNOR2D1 U2647 ( .A1(n2470), .A2(n2441), .Z(n2129) );
  HDNOR2D1 U2648 ( .A1(n2320), .A2(n2755), .Z(n2470) );
  HDOAI211D1 U2649 ( .A1(n2127), .A2(n2443), .B(n2346), .C(n2126), .Z(n2133)
         );
  HDNOR3D1 U2650 ( .A1(n2263), .A2(n2125), .A3(n2826), .Z(n2126) );
  HDNOR2D1 U2651 ( .A1(n2618), .A2(n2819), .Z(n2826) );
  HDINVD1 U2652 ( .A(n2851), .Z(n2263) );
  HDNAN4D1 U2653 ( .A1(n2123), .A2(n2122), .A3(n2121), .A4(n2120), .Z(n2134)
         );
  HDNAN2D1 U2654 ( .A1(n2356), .A2(n2696), .Z(n2120) );
  HDAOI211D1 U2655 ( .A1(n2505), .A2(n2119), .B(n2822), .C(n2118), .Z(n2122)
         );
  HDAOI21D1 U2656 ( .A1(n2117), .A2(n2116), .B(n2929), .Z(n2118) );
  HDAOI211D1 U2657 ( .A1(n2115), .A2(n2158), .B(n2114), .C(n1128), .Z(n2116)
         );
  HDNAN2D1 U2658 ( .A1(n2720), .A2(n679), .Z(n2115) );
  HDNOR4D1 U2659 ( .A1(n2112), .A2(n2724), .A3(n2966), .A4(n2111), .Z(n2117)
         );
  HDAND3D1 U2660 ( .A1(n1383), .A2(n1797), .A3(instruction[8]), .Z(n2966) );
  HDINVD1 U2661 ( .A(n2988), .Z(n1797) );
  HDNAN2D1 U2662 ( .A1(n2100), .A2(n633), .Z(n1383) );
  HDAOI31D1 U2663 ( .A1(n2110), .A2(n1139), .A3(n647), .B(n2927), .Z(n2724) );
  HDAOI21D1 U2664 ( .A1(n2965), .A2(n2109), .B(n2108), .Z(n2112) );
  HDINVD1 U2665 ( .A(n2170), .Z(n2726) );
  HDNOR2D1 U2666 ( .A1(n2107), .A2(n1720), .Z(n2822) );
  HDOAI211D1 U2667 ( .A1(instruction[7]), .A2(n2442), .B(n2104), .C(n2103), 
        .Z(n2105) );
  HDINVD1 U2668 ( .A(n2163), .Z(n2183) );
  HDOAI21D1 U2669 ( .A1(n2685), .A2(n2182), .B(n2099), .Z(n2104) );
  HDNOR2D1 U2670 ( .A1(n2901), .A2(n1811), .Z(n2099) );
  HDNOR2D1 U2671 ( .A1(n2098), .A2(instruction[12]), .Z(n2182) );
  HDINVD1 U2672 ( .A(n2675), .Z(n2685) );
  HDNAN2D1 U2673 ( .A1(n2481), .A2(n2982), .Z(n2442) );
  HDOAI22D1 U2674 ( .A1(instruction[12]), .A2(n2140), .B1(n2417), .B2(
        instruction[15]), .Z(n2106) );
  HDOAI211D1 U2675 ( .A1(n2782), .A2(n2781), .B(n2780), .C(n2779), .Z(
        o_rs1_type[1]) );
  HDNAN2D1 U2676 ( .A1(n2360), .A2(n2784), .Z(n2774) );
  HDNAN2D1 U2677 ( .A1(n2881), .A2(n535), .Z(n2775) );
  HDOAI21M20D1 U2678 ( .A1(n1795), .A2(n2883), .B(n399), .Z(n425) );
  HDOAI22D1 U2679 ( .A1(n388), .A2(n2977), .B1(n1794), .B2(n2902), .Z(n1795)
         );
  HDNOR2D1 U2680 ( .A1(n2805), .A2(n2712), .Z(n1794) );
  HDINVD1 U2681 ( .A(n2771), .Z(n2781) );
  HDNOR2D1 U2682 ( .A1(n2861), .A2(n2766), .Z(n2768) );
  HDNAN2D1 U2683 ( .A1(n1719), .A2(n2778), .Z(n2759) );
  HDNAN2D1 U2684 ( .A1(n2511), .A2(n2520), .Z(n2761) );
  HDNOR4D1 U2685 ( .A1(n2135), .A2(n2094), .A3(n2093), .A4(n2092), .Z(n2095)
         );
  HDNAN4D1 U2686 ( .A1(n2091), .A2(n2090), .A3(n2089), .A4(n2088), .Z(n2092)
         );
  HDINVD1 U2687 ( .A(n2975), .Z(n2989) );
  HDINVD1 U2688 ( .A(n2524), .Z(n2778) );
  HDNOR2D1 U2689 ( .A1(n2866), .A2(n2082), .Z(n2820) );
  HDINVD1 U2690 ( .A(n2907), .Z(n2866) );
  HDOAI211D1 U2691 ( .A1(n2081), .A2(n2640), .B(n2080), .C(n2079), .Z(n2093)
         );
  HDOAI31D1 U2692 ( .A1(n2078), .A2(n2077), .A3(n2076), .B(n2881), .Z(n2079)
         );
  HDOAI211D1 U2693 ( .A1(n2075), .A2(n2987), .B(n2074), .C(n2895), .Z(n2076)
         );
  HDNOR2D1 U2694 ( .A1(n2986), .A2(n2988), .Z(n535) );
  HDNOR2D1 U2695 ( .A1(n2959), .A2(n2974), .Z(n2110) );
  HDINVD1 U2696 ( .A(n2158), .Z(n2415) );
  HDOAI211D1 U2697 ( .A1(n2073), .A2(n2108), .B(n2072), .C(n2159), .Z(n2078)
         );
  HDINVD1 U2698 ( .A(n840), .Z(n885) );
  HDNOR2D1 U2699 ( .A1(n834), .A2(n2755), .Z(n2114) );
  HDINVD1 U2700 ( .A(n2111), .Z(n2072) );
  HDINVD1 U2701 ( .A(n2465), .Z(n2108) );
  HDNOR2D1 U2702 ( .A1(n2068), .A2(n1231), .Z(n2073) );
  HDINVD1 U2703 ( .A(n992), .Z(n2068) );
  HDAOI211D1 U2704 ( .A1(n2288), .A2(instruction[14]), .B(n2885), .C(n2067), 
        .Z(n2080) );
  HDAOI21D1 U2705 ( .A1(n2359), .A2(n2798), .B(n2066), .Z(n2067) );
  HDNOR2D1 U2706 ( .A1(n2064), .A2(instruction[12]), .Z(n2065) );
  HDNAN2D1 U2707 ( .A1(instruction[7]), .A2(instruction[5]), .Z(n1811) );
  HDINVD1 U2708 ( .A(n2725), .Z(n2100) );
  HDNOR2D1 U2709 ( .A1(n2851), .A2(n2982), .Z(n2885) );
  HDNOR2D1 U2710 ( .A1(n1644), .A2(instruction[6]), .Z(n2063) );
  HDINVD1 U2711 ( .A(n2925), .Z(n2062) );
  HDINVD1 U2712 ( .A(n2417), .Z(n2288) );
  HDNOR2D1 U2713 ( .A1(n2799), .A2(n2319), .Z(n2058) );
  HDNOR2D1 U2714 ( .A1(n2982), .A2(instruction[7]), .Z(n2319) );
  HDNAN2D1 U2715 ( .A1(n2980), .A2(instruction[13]), .Z(n2060) );
  HDOAI211D1 U2716 ( .A1(n2320), .A2(n2853), .B(n2051), .C(n2050), .Z(n2094)
         );
  HDNOR2D1 U2717 ( .A1(n2767), .A2(instruction[28]), .Z(n2048) );
  HDINVD1 U2718 ( .A(n2140), .Z(n2047) );
  HDINVD1 U2719 ( .A(n415), .Z(n2853) );
  HDNAN4D1 U2720 ( .A1(n2045), .A2(n2044), .A3(n2043), .A4(n2343), .Z(n2135)
         );
  HDNOR2D1 U2721 ( .A1(n2280), .A2(n2042), .Z(n2343) );
  HDAOI211D1 U2722 ( .A1(n2171), .A2(n2308), .B(n2039), .C(n2038), .Z(n2045)
         );
  HDNOR4D1 U2723 ( .A1(n2037), .A2(n2036), .A3(n2453), .A4(n2035), .Z(n2096)
         );
  HDNOR2D1 U2724 ( .A1(n2236), .A2(n2951), .Z(n2234) );
  HDNOR2D1 U2725 ( .A1(instruction[23]), .A2(instruction[22]), .Z(n2453) );
  HDNOR4D1 U2726 ( .A1(n2031), .A2(n1697), .A3(n2325), .A4(n2148), .Z(n2033)
         );
  HDINVD1 U2727 ( .A(n2029), .Z(n2236) );
  HDOAI211D1 U2728 ( .A1(instruction[28]), .A2(n2321), .B(n2550), .C(n2209), 
        .Z(n2326) );
  HDNOR4D1 U2729 ( .A1(n2589), .A2(n1697), .A3(n2146), .A4(n2219), .Z(n2209)
         );
  HDNOR4D1 U2730 ( .A1(n2028), .A2(n2027), .A3(n2406), .A4(n2026), .Z(n2097)
         );
  HDNAN2D1 U2731 ( .A1(n1867), .A2(n1866), .Z(n2025) );
  HDNOR4D1 U2732 ( .A1(n1796), .A2(n387), .A3(instruction[13]), .A4(n2980), 
        .Z(n1866) );
  HDAOI211D1 U2733 ( .A1(n1685), .A2(n1863), .B(n2441), .C(n1862), .Z(n2023)
         );
  HDINVD1 U2734 ( .A(n2407), .Z(n2271) );
  HDNOR2D1 U2735 ( .A1(n1861), .A2(n2199), .Z(n2441) );
  HDINVD1 U2736 ( .A(n2138), .Z(n2024) );
  HDNAN2D1 U2737 ( .A1(n2256), .A2(n2257), .Z(n2346) );
  HDOR4D1 U2738 ( .A1(n1668), .A2(n1970), .A3(n1971), .A4(n1728), .Z(
        o_m_imm[31]) );
  HDOAI211D1 U2739 ( .A1(n2868), .A2(n2374), .B(n1968), .C(n1967), .Z(n1668)
         );
  HDNAN2D1 U2740 ( .A1(n2497), .A2(instruction[29]), .Z(n1968) );
  HDNAN2M1D1 U2741 ( .A1(n1664), .A2(n1656), .Z(n1654) );
  HDOAI21D1 U2742 ( .A1(n2740), .A2(n2977), .B(n2804), .Z(n2933) );
  HDNAN2D1 U2743 ( .A1(n2800), .A2(n2902), .Z(n2804) );
  HDOAI22M10D1 U2744 ( .A1(n1663), .A2(n2930), .B1(n1658), .B2(n2929), .Z(
        n1657) );
  HDAND2D1 U2745 ( .A1(n1641), .A2(n1646), .Z(n2719) );
  HDAND4D1 U2746 ( .A1(n1642), .A2(n2785), .A3(n2924), .A4(n1643), .Z(n1646)
         );
  HDOR2D1 U2747 ( .A1(n2988), .A2(instruction[8]), .Z(n1643) );
  HDNOR2D1 U2748 ( .A1(n2979), .A2(n930), .Z(n2274) );
  HDNOR2D1 U2749 ( .A1(n2982), .A2(n2981), .Z(n1230) );
  HDOAI21D1 U2750 ( .A1(n2927), .A2(n2720), .B(n679), .Z(n1620) );
  HDNOR2D1 U2751 ( .A1(n2718), .A2(n2784), .Z(n2722) );
  HDNOR2D1 U2752 ( .A1(n2465), .A2(n2787), .Z(n2718) );
  HDINVD1 U2753 ( .A(n1796), .Z(n2787) );
  HDOAI211D1 U2754 ( .A1(n2979), .A2(n2980), .B(n681), .C(n2982), .Z(n674) );
  HDINVD1 U2755 ( .A(n595), .Z(n2974) );
  HDAND2D1 U2756 ( .A1(n2113), .A2(n2980), .Z(n2975) );
  HDNAN2D1 U2757 ( .A1(n2742), .A2(n2741), .Z(n2922) );
  HDAND2D1 U2758 ( .A1(n1807), .A2(n2101), .Z(n2098) );
  HDAND2D1 U2759 ( .A1(n595), .A2(n2727), .Z(n2923) );
  HDNOR4D1 U2760 ( .A1(n1652), .A2(n1662), .A3(n2920), .A4(n2921), .Z(n1655)
         );
  HDINVD1 U2761 ( .A(n2749), .Z(n2917) );
  HDINVD1 U2762 ( .A(n2186), .Z(n2918) );
  HDOAI211D1 U2763 ( .A1(n2016), .A2(n2934), .B(n2015), .C(n2014), .Z(
        o_m_branch_type[1]) );
  HDOAI211D1 U2764 ( .A1(instruction[29]), .A2(n2216), .B(n2012), .C(n2011), 
        .Z(n2013) );
  HDOR4D1 U2765 ( .A1(n1976), .A2(o_rs2_2_), .A3(o_rs2_4_), .A4(n1975), .Z(
        n2011) );
  HDNAN4D1 U2766 ( .A1(n2175), .A2(instruction[13]), .A3(n1443), .A4(o_rs2_3_), 
        .Z(n1975) );
  HDINVD1 U2767 ( .A(n2128), .Z(n2012) );
  HDINVD1 U2768 ( .A(n2010), .Z(n2216) );
  HDINVD1 U2769 ( .A(n2339), .Z(n2380) );
  HDNAN4D1 U2770 ( .A1(n2534), .A2(n2637), .A3(n2576), .A4(n2840), .Z(
        o_rs4_valid) );
  HDINVD1 U2771 ( .A(o_m_flags[2]), .Z(n2576) );
  HDINVD1 U2772 ( .A(n2583), .Z(n1867) );
  HDNAN2D1 U2773 ( .A1(n2082), .A2(n2696), .Z(n2583) );
  HDNAN3D1 U2774 ( .A1(n2577), .A2(n1834), .A3(n2450), .Z(n1836) );
  HDNOR3D1 U2775 ( .A1(n1696), .A2(n1833), .A3(n2749), .Z(n1834) );
  HDINVD1 U2776 ( .A(n2520), .Z(n1833) );
  HDINVD1 U2777 ( .A(n2818), .Z(n1696) );
  HDINVD1 U2778 ( .A(n2762), .Z(n2818) );
  HDAND4D1 U2779 ( .A1(n2764), .A2(n2511), .A3(n1747), .A4(n2676), .Z(n2577)
         );
  HDNOR2D1 U2780 ( .A1(n2187), .A2(n2408), .Z(n1747) );
  HDINVD1 U2781 ( .A(n2872), .Z(n2187) );
  HDNOR2D1 U2782 ( .A1(n2634), .A2(n2572), .Z(n2529) );
  HDNAN2D1 U2783 ( .A1(n1853), .A2(n2673), .Z(n2572) );
  HDINVD1 U2784 ( .A(n2924), .Z(n2905) );
  HDOR2D1 U2785 ( .A1(n387), .A2(n1644), .Z(n2924) );
  HDINVD1 U2786 ( .A(n1229), .Z(n1644) );
  HDNOR2D1 U2787 ( .A1(n2610), .A2(n2528), .Z(n2571) );
  HDINVD1 U2788 ( .A(n2730), .Z(n2610) );
  HDINVD1 U2789 ( .A(n2085), .Z(n1760) );
  HDNOR4D1 U2790 ( .A1(n2567), .A2(n2547), .A3(n2590), .A4(n2527), .Z(n2531)
         );
  HDNAN2D1 U2791 ( .A1(n2628), .A2(n2604), .Z(n2527) );
  HDINVD1 U2792 ( .A(n2609), .Z(n2547) );
  HDAND2D1 U2793 ( .A1(n2425), .A2(n2308), .Z(n2860) );
  HDAND2D1 U2794 ( .A1(n2323), .A2(n2258), .Z(n2308) );
  HDNAN3D1 U2795 ( .A1(n1686), .A2(n2175), .A3(n2812), .Z(n2425) );
  HDINVD1 U2796 ( .A(n2285), .Z(n2175) );
  HDINVD1 U2797 ( .A(n2054), .Z(n2561) );
  HDOAI211D1 U2798 ( .A1(n2054), .A2(n2810), .B(n2615), .C(n2633), .Z(n2545)
         );
  HDNAN4D1 U2799 ( .A1(n2558), .A2(n2630), .A3(n2562), .A4(n2625), .Z(n1851)
         );
  HDNOR2D1 U2800 ( .A1(n2052), .A2(n2797), .Z(n2542) );
  HDNAN2D1 U2801 ( .A1(n2812), .A2(instruction[17]), .Z(n2052) );
  HDNOR2D1 U2802 ( .A1(n2540), .A2(n2535), .Z(n2562) );
  HDAND3D1 U2803 ( .A1(n2771), .A2(n2310), .A3(instruction[14]), .Z(n2535) );
  HDNOR2D1 U2804 ( .A1(n2556), .A2(n2559), .Z(n2630) );
  HDNOR2D1 U2805 ( .A1(n1848), .A2(n2160), .Z(n2559) );
  HDNAN2D1 U2806 ( .A1(instruction[15]), .A2(instruction[16]), .Z(n2160) );
  HDNOR2D1 U2807 ( .A1(n2281), .A2(n1847), .Z(n2556) );
  HDNAN2D1 U2808 ( .A1(n1846), .A2(instruction[15]), .Z(n2281) );
  HDAOI21D1 U2809 ( .A1(n2287), .A2(n2812), .B(n2599), .Z(n2558) );
  HDNOR2D1 U2810 ( .A1(n2284), .A2(instruction[18]), .Z(n2599) );
  HDNAN3D1 U2811 ( .A1(n2537), .A2(instruction[14]), .A3(instruction[16]), .Z(
        n2284) );
  HDNAN2D1 U2812 ( .A1(n2053), .A2(n2285), .Z(n1841) );
  HDNAN3D1 U2813 ( .A1(n2317), .A2(instruction[16]), .A3(instruction[17]), .Z(
        n2285) );
  HDAND2D1 U2814 ( .A1(instruction[14]), .A2(instruction[15]), .Z(n2317) );
  HDOAI211D1 U2815 ( .A1(n2543), .A2(n2310), .B(n1840), .C(n2811), .Z(n2053)
         );
  HDINVD1 U2816 ( .A(n1846), .Z(n1848) );
  HDNAN2D1 U2817 ( .A1(n2287), .A2(instruction[18]), .Z(n1844) );
  HDNAN2D1 U2818 ( .A1(n2538), .A2(n2626), .Z(n2287) );
  HDNAN2D1 U2819 ( .A1(n1846), .A2(n2310), .Z(n2538) );
  HDNAN2D1 U2820 ( .A1(instruction[14]), .A2(instruction[17]), .Z(n1845) );
  HDINVD1 U2821 ( .A(n1847), .Z(n2536) );
  HDOR2D1 U2822 ( .A1(instruction[18]), .A2(instruction[16]), .Z(n1847) );
  HDNAN2D1 U2823 ( .A1(n2537), .A2(n1840), .Z(n2054) );
  HDAND2D1 U2824 ( .A1(instruction[14]), .A2(instruction[18]), .Z(n1840) );
  HDOAI211D1 U2825 ( .A1(n1936), .A2(n1947), .B(n1925), .C(n1924), .Z(
        o_m_imm[11]) );
  HDAOI211D1 U2826 ( .A1(n1923), .A2(instruction[11]), .B(n1608), .C(n1728), 
        .Z(n1924) );
  HDNAN2D1 U2827 ( .A1(n2876), .A2(o_rs2_1_), .Z(n1925) );
  HDOAI211D1 U2828 ( .A1(n2868), .A2(n2064), .B(n1674), .C(n1955), .Z(
        o_m_imm[21]) );
  HDNAN2D1 U2829 ( .A1(n1954), .A2(instruction[19]), .Z(n1674) );
  HDOAI211D1 U2830 ( .A1(n2868), .A2(n2399), .B(n1675), .C(n1955), .Z(
        o_m_imm[22]) );
  HDNOR2D4 U2831 ( .A1(n1728), .A2(n1971), .Z(n1964) );
  HDNAN3D1 U2832 ( .A1(n2941), .A2(instruction[18]), .A3(n2217), .Z(n1952) );
  HDNAN2D1 U2833 ( .A1(n2770), .A2(instruction[21]), .Z(n1953) );
  HDAOI211D1 U2834 ( .A1(n1686), .A2(n1731), .B(n1888), .C(n2257), .Z(n1889)
         );
  HDOR2D1 U2835 ( .A1(n1909), .A2(n1911), .Z(n1617) );
  HDNAN3D1 U2836 ( .A1(n2738), .A2(n2939), .A3(instruction[13]), .Z(n1911) );
  HDOAI22D1 U2837 ( .A1(n2640), .A2(n2978), .B1(n2798), .B2(n1947), .Z(n1909)
         );
  HDAOI211D1 U2838 ( .A1(n2597), .A2(n2506), .B(n2408), .C(n1800), .Z(n1801)
         );
  HDINVD1 U2839 ( .A(n2202), .Z(n2087) );
  HDAND4D1 U2840 ( .A1(n1669), .A2(n1825), .A3(n2525), .A4(n1670), .Z(n1672)
         );
  HDINVD1 U2841 ( .A(n2883), .Z(n1670) );
  HDINVD1 U2842 ( .A(n2309), .Z(n2192) );
  HDNAN2D1 U2843 ( .A1(n2524), .A2(n2659), .Z(n1863) );
  HDNOR4D1 U2844 ( .A1(n1877), .A2(n1821), .A3(n1820), .A4(n1671), .Z(n1669)
         );
  HDNAN2D1 U2845 ( .A1(n1824), .A2(n2733), .Z(n1671) );
  HDINVD1 U2846 ( .A(n2644), .Z(n1824) );
  HDNAN3D1 U2847 ( .A1(n2767), .A2(n2732), .A3(n2128), .Z(n1820) );
  HDNAN2D1 U2848 ( .A1(n2640), .A2(n2690), .Z(n1877) );
  HDNAN4D1 U2849 ( .A1(n2763), .A2(n2511), .A3(n2458), .A4(n1886), .Z(n1890)
         );
  HDNOR2D1 U2850 ( .A1(n2870), .A2(n2478), .Z(n1886) );
  HDNAN2D1 U2851 ( .A1(n1596), .A2(n2889), .Z(n1883) );
  HDNAN4D1 U2852 ( .A1(n2383), .A2(n1882), .A3(n2459), .A4(n1881), .Z(n1884)
         );
  HDINVD1 U2853 ( .A(n2406), .Z(n1881) );
  HDNOR2D1 U2854 ( .A1(n2921), .A2(n2408), .Z(n1882) );
  HDINVD1 U2855 ( .A(n2673), .Z(n2921) );
  HDOR4D1 U2856 ( .A1(n2648), .A2(n1919), .A3(n2494), .A4(n1666), .Z(n1667) );
  HDINVD1 U2857 ( .A(n2504), .Z(n1771) );
  HDNAN2D1 U2858 ( .A1(n1954), .A2(instruction[20]), .Z(n1675) );
  HDBUFD2 U2859 ( .A(n2777), .Z(n1685) );
  HDOAI211D1 U2860 ( .A1(n2953), .A2(n2946), .B(n1600), .C(n2945), .Z(o_rd[1])
         );
  HDNOR2D1 U2861 ( .A1(n2916), .A2(n1732), .Z(n2947) );
  HDOAI211D1 U2862 ( .A1(n2940), .A2(n2939), .B(n2938), .C(n2937), .Z(n2942)
         );
  HDINVD1 U2863 ( .A(n2936), .Z(n2937) );
  HDNAN2D1 U2864 ( .A1(n1865), .A2(n1888), .Z(n2733) );
  HDAND2D1 U2865 ( .A1(n2817), .A2(n2128), .Z(n2730) );
  HDNAN4D1 U2866 ( .A1(n2919), .A2(n2863), .A3(n2508), .A4(n2507), .Z(n2737)
         );
  HDNOR2D1 U2867 ( .A1(n2506), .A2(n2505), .Z(n2507) );
  HDNOR2D1 U2868 ( .A1(n2679), .A2(instruction[21]), .Z(n1819) );
  HDNOR2D1 U2869 ( .A1(n2198), .A2(n2243), .Z(n2266) );
  HDNAN3D1 U2870 ( .A1(n2437), .A2(n2655), .A3(n2872), .Z(n2504) );
  HDOR2D1 U2871 ( .A1(n2578), .A2(n1706), .Z(n2872) );
  HDINVD1 U2872 ( .A(n2935), .Z(n2940) );
  HDOR2D1 U2873 ( .A1(o_m_branch_type[3]), .A2(n1711), .Z(o_m_type[1]) );
  HDOR3D1 U2874 ( .A1(n2533), .A2(o_m_branch_type[2]), .A3(n2526), .Z(n1711)
         );
  HDNOR2D1 U2875 ( .A1(n2845), .A2(n2200), .Z(n2525) );
  HDNOR2D1 U2876 ( .A1(n1869), .A2(n1868), .Z(n2200) );
  HDNOR3D1 U2877 ( .A1(n2523), .A2(n2522), .A3(n2869), .Z(n2867) );
  HDNAN2D1 U2878 ( .A1(n2375), .A2(n1865), .Z(n2582) );
  HDNOR3D1 U2879 ( .A1(n2408), .A2(n2407), .A3(n2406), .Z(n2521) );
  HDNOR2D1 U2880 ( .A1(n1835), .A2(n1704), .Z(n2407) );
  HDNAN3D1 U2881 ( .A1(n2477), .A2(n2476), .A3(n2475), .Z(n2523) );
  HDAOI211D1 U2882 ( .A1(n2375), .A2(n2374), .B(n2373), .C(n2372), .Z(n2476)
         );
  HDNAN2D1 U2883 ( .A1(n2374), .A2(instruction[20]), .Z(n1706) );
  HDOAI21D1 U2884 ( .A1(n1981), .A2(n2323), .B(n2941), .Z(n1937) );
  HDNOR3D1 U2885 ( .A1(o_m_type[2]), .A2(n2497), .A3(n2496), .Z(n1683) );
  HDOAI211D1 U2886 ( .A1(n2601), .A2(n1732), .B(n2753), .C(n1977), .Z(n2496)
         );
  HDNAN2D1 U2887 ( .A1(n2941), .A2(n2217), .Z(n1977) );
  HDNOR2D1 U2888 ( .A1(n1951), .A2(instruction[23]), .Z(n2217) );
  HDINVD1 U2889 ( .A(n2770), .Z(n2753) );
  HDNAN2D2 U2890 ( .A1(n1951), .A2(instruction[23]), .Z(n2377) );
  HDNAN2D1 U2891 ( .A1(n2491), .A2(n2490), .Z(n1684) );
  HDNOR2D1 U2892 ( .A1(n2481), .A2(n2865), .Z(n2490) );
  HDINVD1 U2893 ( .A(n1161), .Z(n2101) );
  HDNAN2D1 U2894 ( .A1(n2467), .A2(n2881), .Z(n2491) );
  HDOAI211D1 U2895 ( .A1(n1405), .A2(n2987), .B(n2927), .C(n2466), .Z(n2467)
         );
  HDOR2D1 U2896 ( .A1(n388), .A2(n2979), .Z(n992) );
  HDINVD1 U2897 ( .A(n591), .Z(n2983) );
  HDOR2D4 U2898 ( .A1(instruction[30]), .A2(instruction[31]), .Z(n2934) );
  HDNAN2D1 U2899 ( .A1(n2510), .A2(n2265), .Z(n2907) );
  HDMUX2D1 U2900 ( .A0(n1679), .A1(n1680), .SL(n2570), .Z(n2515) );
  HDINVD1 U2901 ( .A(n2244), .Z(n2324) );
  HDNOR2D1 U2902 ( .A1(n2148), .A2(n2006), .Z(n2246) );
  HDINVD1 U2903 ( .A(n2617), .Z(n1719) );
  HDNOR2D1 U2904 ( .A1(n1678), .A2(n2589), .Z(n1677) );
  HDOR2D1 U2905 ( .A1(n1999), .A2(n2746), .Z(n1676) );
  HDNOR2D1 U2906 ( .A1(n1697), .A2(n2000), .Z(n2214) );
  HDOAI211D1 U2907 ( .A1(n1999), .A2(n1998), .B(n1997), .C(n1996), .Z(n2003)
         );
  HDINVD1 U2908 ( .A(n1994), .Z(n1997) );
  HDNAN2M1D1 U2909 ( .A1(n1727), .A2(n1993), .Z(n2624) );
  HDAOI211D1 U2910 ( .A1(n2009), .A2(instruction[5]), .B(n2000), .C(n2006), 
        .Z(n1993) );
  HDINVD1 U2911 ( .A(n1989), .Z(n2000) );
  HDAND2D1 U2912 ( .A1(n2147), .A2(n2948), .Z(n2589) );
  HDNOR2D1 U2913 ( .A1(n1689), .A2(instruction[28]), .Z(n2147) );
  HDNOR2D1 U2914 ( .A1(n2944), .A2(n2242), .Z(n2146) );
  HDNAN2D1 U2915 ( .A1(n1995), .A2(n2617), .Z(n1987) );
  HDNAN2D1 U2916 ( .A1(n1985), .A2(n1984), .Z(n2244) );
  HDOAI211D1 U2917 ( .A1(n1983), .A2(n2952), .B(n1989), .C(n1982), .Z(n1988)
         );
  HDAO21M20D1 U2918 ( .A1(n2212), .A2(n2325), .B(instruction[29]), .Z(n1982)
         );
  HDNAN2D1 U2919 ( .A1(n1984), .A2(n2210), .Z(n1989) );
  HDINVD1 U2920 ( .A(n2943), .Z(n1984) );
  HDNOR4D1 U2921 ( .A1(n2030), .A2(n2339), .A3(n2231), .A4(n2001), .Z(n1983)
         );
  HDINVD1 U2922 ( .A(n2379), .Z(n2162) );
  HDNOR2D1 U2923 ( .A1(n1992), .A2(n2031), .Z(n2007) );
  HDINVD1 U2924 ( .A(n1991), .Z(n2031) );
  HDNOR2D1 U2925 ( .A1(n2219), .A2(n2010), .Z(n1991) );
  HDNOR2D1 U2926 ( .A1(n1689), .A2(n1986), .Z(n2010) );
  HDNOR2D1 U2927 ( .A1(n2242), .A2(n2379), .Z(n2219) );
  HDOR2D1 U2928 ( .A1(instruction[26]), .A2(instruction[25]), .Z(n2379) );
  HDINVD1 U2929 ( .A(n2325), .Z(n2233) );
  HDNOR2D1 U2930 ( .A1(n2714), .A2(n2939), .Z(n2758) );
  HDNOR2D1 U2931 ( .A1(n2935), .A2(instruction[8]), .Z(n2712) );
  HDINVD1 U2932 ( .A(n2059), .Z(n2805) );
  HDNOR4D1 U2933 ( .A1(n2064), .A2(n1947), .A3(instruction[13]), .A4(
        instruction[10]), .Z(n1761) );
  HDOAI211D1 U2934 ( .A1(n2709), .A2(n2755), .B(n2708), .C(n2707), .Z(n2710)
         );
  HDAOI22D1 U2935 ( .A1(n2899), .A2(n409), .B1(n1763), .B2(n2158), .Z(n2707)
         );
  HDNAN2D1 U2936 ( .A1(n2170), .A2(n679), .Z(n1763) );
  HDNAN2D1 U2937 ( .A1(n2979), .A2(n840), .Z(n679) );
  HDNOR2D1 U2938 ( .A1(n2982), .A2(n2981), .Z(n1702) );
  HDOR2D1 U2939 ( .A1(n633), .A2(instruction[8]), .Z(n2170) );
  HDOR2D1 U2940 ( .A1(n387), .A2(n1738), .Z(n595) );
  HDNAN2M1D1 U2941 ( .A1(instruction[8]), .A2(instruction[7]), .Z(n1738) );
  HDNAN2D1 U2942 ( .A1(n2927), .A2(n2988), .Z(n2706) );
  HDNOR2D1 U2943 ( .A1(n416), .A2(n2465), .Z(n2709) );
  HDNOR2D1 U2944 ( .A1(n2086), .A2(instruction[12]), .Z(n2465) );
  HDNAN2D1 U2945 ( .A1(n2978), .A2(instruction[11]), .Z(n1807) );
  HDNAN2D1 U2946 ( .A1(n835), .A2(n834), .Z(n416) );
  HDNAN2D1 U2947 ( .A1(n2928), .A2(n1229), .Z(n834) );
  HDNOR2D1 U2948 ( .A1(instruction[8]), .A2(instruction[7]), .Z(n1229) );
  HDNOR3D1 U2949 ( .A1(n2675), .A2(instruction[10]), .A3(n1947), .Z(n2928) );
  HDNAN2D1 U2950 ( .A1(instruction[11]), .A2(instruction[12]), .Z(n2675) );
  HDOR2D1 U2951 ( .A1(n2399), .A2(instruction[9]), .Z(n1708) );
  HDNAN2D1 U2952 ( .A1(n2978), .A2(instruction[11]), .Z(n1707) );
  HDAND2D1 U2953 ( .A1(n2713), .A2(instruction[8]), .Z(n2959) );
  HDNOR2D1 U2954 ( .A1(o_rs2_4_), .A2(o_rs2_3_), .Z(n2716) );
  HDNOR2D1 U2955 ( .A1(n2510), .A2(n2039), .Z(n2520) );
  HDINVD1 U2956 ( .A(n2019), .Z(n2039) );
  HDOAI211D1 U2957 ( .A1(instruction[19]), .A2(n2199), .B(n1860), .C(n1778), 
        .Z(n1779) );
  HDINVD1 U2958 ( .A(n2422), .Z(n2348) );
  HDNAN2D1 U2959 ( .A1(n2257), .A2(n1865), .Z(n2422) );
  HDNAN2D1 U2960 ( .A1(n1688), .A2(n2578), .Z(n2145) );
  HDINVD1 U2961 ( .A(n2257), .Z(n2199) );
  HDNAN4D1 U2962 ( .A1(n1776), .A2(n2674), .A3(n2889), .A4(n2382), .Z(n1919)
         );
  HDNAN3D1 U2963 ( .A1(n2265), .A2(n2018), .A3(n1731), .Z(n2495) );
  HDINVD1 U2964 ( .A(n2475), .Z(n2892) );
  HDNAN2D1 U2965 ( .A1(n2511), .A2(n2383), .Z(n1780) );
  HDNAN3D1 U2966 ( .A1(n1775), .A2(n2641), .A3(n2083), .Z(n1781) );
  HDAND3D1 U2967 ( .A1(n2330), .A2(n2361), .A3(n2673), .Z(n2083) );
  HDNOR2D1 U2968 ( .A1(n2125), .A2(n2040), .Z(n2641) );
  HDINVD1 U2969 ( .A(n2464), .Z(n2125) );
  HDINVD1 U2970 ( .A(n2136), .Z(n1775) );
  HDNAN3D1 U2971 ( .A1(n2874), .A2(n2435), .A3(n1853), .Z(n2136) );
  HDINVD1 U2972 ( .A(n2760), .Z(n2874) );
  HDOAI21D1 U2973 ( .A1(n2703), .A2(n2861), .B(n1609), .Z(n2704) );
  HDAND2D4 U2974 ( .A1(n1892), .A2(instruction[31]), .Z(n1609) );
  HDNOR2D1 U2975 ( .A1(n2979), .A2(instruction[7]), .Z(n1395) );
  HDINVBD4 U2976 ( .A(instruction[8]), .Z(n2979) );
  HDAOI21D1 U2977 ( .A1(n2769), .A2(n2702), .B(instruction[13]), .Z(n2703) );
  HDNOR3D1 U2978 ( .A1(n2858), .A2(n2766), .A3(n2356), .Z(n2702) );
  HDNOR3D1 U2979 ( .A1(n2658), .A2(n1773), .A3(n1812), .Z(n2766) );
  HDINVD1 U2980 ( .A(n1888), .Z(n1773) );
  HDNAN3D1 U2981 ( .A1(n2471), .A2(n2798), .A3(n2640), .Z(n2858) );
  HDINVBD4 U2982 ( .A(n2795), .Z(n2798) );
  HDAND2D1 U2983 ( .A1(n2189), .A2(n2323), .Z(n2506) );
  HDAND2D1 U2984 ( .A1(n2124), .A2(n2809), .Z(n2444) );
  HDNOR2D1 U2985 ( .A1(instruction[14]), .A2(instruction[16]), .Z(n2124) );
  HDINVD1 U2986 ( .A(n2528), .Z(n2699) );
  HDNAN2D1 U2987 ( .A1(n2383), .A2(n2382), .Z(n2528) );
  HDNAN2M1D1 U2988 ( .A1(n2578), .A2(n2500), .Z(n2382) );
  HDAND3D1 U2989 ( .A1(n2259), .A2(n2202), .A3(n2472), .Z(n2383) );
  HDOR2D1 U2990 ( .A1(n2327), .A2(n1713), .Z(n2472) );
  HDNAN2D1 U2991 ( .A1(n2256), .A2(n1822), .Z(n2202) );
  HDNAN2D1 U2992 ( .A1(n1873), .A2(n2500), .Z(n2259) );
  HDINVD1 U2993 ( .A(n2698), .Z(n2700) );
  HDNAN2D1 U2994 ( .A1(n2601), .A2(n2128), .Z(n2698) );
  HDAND2D1 U2995 ( .A1(n1770), .A2(n1731), .Z(n2460) );
  HDAND2D1 U2996 ( .A1(n1749), .A2(n2374), .Z(n1770) );
  HDNAN2D1 U2997 ( .A1(instruction[20]), .A2(instruction[19]), .Z(n1749) );
  HDINVD1 U2998 ( .A(n2459), .Z(n2461) );
  HDNAN2D1 U2999 ( .A1(n1731), .A2(n1712), .Z(n2493) );
  HDNAN2D4 U3000 ( .A1(n1823), .A2(n1731), .Z(n2673) );
  HDNOR2D2 U3001 ( .A1(instruction[23]), .A2(instruction[24]), .Z(n1777) );
  HDOR2D1 U3002 ( .A1(n1688), .A2(n1713), .Z(n2361) );
  HDNOR2D1 U3003 ( .A1(n1831), .A2(n1687), .Z(n2038) );
  HDINVD1 U3004 ( .A(n1774), .Z(n1712) );
  HDNAN2D2 U3005 ( .A1(instruction[21]), .A2(instruction[20]), .Z(n1774) );
  HDOR2D1 U3006 ( .A1(n1753), .A2(n1687), .Z(n2330) );
  HDNOR3D4 U3007 ( .A1(instruction[19]), .A2(instruction[21]), .A3(
        instruction[20]), .Z(n2258) );
  HDNOR2D1 U3008 ( .A1(n2338), .A2(n1868), .Z(n2042) );
  HDNAN3D2 U3009 ( .A1(n1746), .A2(n2374), .A3(instruction[20]), .Z(n1868) );
  HDNOR3D4 U3010 ( .A1(n1746), .A2(instruction[21]), .A3(instruction[20]), .Z(
        n2501) );
  HDOR2D4 U3011 ( .A1(n1740), .A2(instruction[22]), .Z(n2243) );
  HDAND2DL U3012 ( .A1(n1870), .A2(n1599), .Z(o_m_access_size[4]) );
  HDOAI21M20DL U3013 ( .A1(n2830), .A2(n2849), .B(n2829), .Z(o_rd2_type[1]) );
  HDOAI21M20DL U3014 ( .A1(N5188), .A2(n2849), .B(n2847), .Z(o_rd2[4]) );
  HDOAI21M20DL U3015 ( .A1(n2479), .A2(n1609), .B(n2489), .Z(o_m_futype[0]) );
  HDNAN2DL U3016 ( .A1(n2789), .A2(n2727), .Z(n2728) );
  HDOAI21M20DL U3017 ( .A1(n2973), .A2(instruction[8]), .B(n2100), .Z(n1764)
         );
  HDAOI22DL U3018 ( .A1(n2492), .A2(n2219), .B1(n2218), .B2(n2217), .Z(n2220)
         );
  HDOAI21M20DL U3019 ( .A1(n2214), .A2(n2321), .B(n2323), .Z(n2221) );
  HDOAI21M20DL U3020 ( .A1(n2320), .A2(n2177), .B(n2982), .Z(n2178) );
  HDOAI21M20DL U3021 ( .A1(n1084), .A2(n2176), .B(n2481), .Z(n2177) );
  HDEXNOR2DL U3022 ( .A1(instruction[14]), .A2(instruction[15]), .Z(n2166) );
  HDAOI22DL U3023 ( .A1(n1888), .A2(n2941), .B1(n2770), .B2(instruction[28]), 
        .Z(n1827) );
  HDAOI211DL U3024 ( .A1(n1630), .A2(n2322), .B(n2453), .C(n1631), .Z(n1628)
         );
  HDAND4DL U3025 ( .A1(n2426), .A2(n2309), .A3(n2418), .A4(n1824), .Z(n1622)
         );
  HDOAI21M20DL U3026 ( .A1(n2717), .A2(n2716), .B(n2715), .Z(o_rs2_type[1]) );
  HDMUXB2DL U3027 ( .A0(n2797), .A1(n2796), .SL(n1609), .Z(o_rs1[0]) );
  HDMUXB2DL U3028 ( .A0(n633), .A1(n885), .SL(n2352), .Z(n2354) );
  HDOAI21M20DL U3029 ( .A1(n1794), .A2(n2060), .B(n2883), .Z(n1762) );
  HDOAI21M20DL U3030 ( .A1(n1787), .A2(instruction[14]), .B(n2901), .Z(n1788)
         );
  HDNAN3DL U3031 ( .A1(n1716), .A2(n1964), .A3(n1961), .Z(o_m_imm[28]) );
  HDNAN3DL U3032 ( .A1(n1965), .A2(n1964), .A3(n1962), .Z(o_m_imm[29]) );
  HDNAN3DL U3033 ( .A1(n1965), .A2(n1964), .A3(n1963), .Z(o_m_imm[30]) );
  HDNAN2DL U3034 ( .A1(n2257), .A2(n2189), .Z(n2349) );
  HDOAI21M20DL U3035 ( .A1(n2234), .A2(n2233), .B(n2323), .Z(n2239) );
  HDOAI21M20DL U3036 ( .A1(n2800), .A2(n2797), .B(n2663), .Z(n2665) );
  HDNAN2DL U3037 ( .A1(n2266), .A2(n2265), .Z(n2398) );
  HDAOI21M20DL U3038 ( .A1(n2393), .A2(n2392), .B(n2391), .Z(n2395) );
  HDOAI21DL U3039 ( .A1(n2971), .A2(n1231), .B(n2865), .Z(n2089) );
  HDAOI21M20DL U3040 ( .A1(n834), .A2(n1137), .B(n535), .Z(n2074) );
  HDMUXB2DL U3041 ( .A0(instruction[12]), .A1(n2065), .SL(n2978), .Z(n2066) );
  HDAOI21M20DL U3042 ( .A1(n2310), .A2(instruction[14]), .B(n2052), .Z(n2057)
         );
  HDMUXB2DL U3043 ( .A0(n2047), .A1(n2748), .SL(n2399), .Z(n2051) );
  HDEXOR2DL U3044 ( .A1(instruction[28]), .A2(instruction[25]), .Z(n2034) );
  HDMUXB2DL U3045 ( .A0(n1161), .A1(n1544), .SL(instruction[9]), .Z(n2741) );
  HDOAI21M20DL U3046 ( .A1(n2944), .A2(n2943), .B(n2947), .Z(n2945) );
  HDINVD1 U3047 ( .A(o_rs2_3_), .Z(n1998) );
  HDMUXB2DL U3048 ( .A0(n2799), .A1(n2319), .SL(n2352), .Z(n1640) );
  HDNAN3DL U3049 ( .A1(n2731), .A2(n2511), .A3(n2733), .Z(n1652) );
  HDAO211DL U3050 ( .A1(n2925), .A2(n2924), .B(n2923), .C(n2922), .Z(n1663) );
  HDTIELO U3051 ( .Z(n_Logic0_) );
  HDINVD1 U3052 ( .A(instruction[26]), .Z(n2946) );
  HDAOI22DL U3053 ( .A1(n2258), .A2(n2257), .B1(n2375), .B2(n2256), .Z(n2260)
         );
  HDAOI21M20DL U3054 ( .A1(n2326), .A2(n2236), .B(n1688), .Z(n2037) );
  HDAOI21DL U3055 ( .A1(n2883), .A2(n388), .B(n2739), .Z(n2740) );
  HDAOI21M20DL U3056 ( .A1(n2237), .A2(n2210), .B(n2243), .Z(n2225) );
  HDAOI21M20DL U3057 ( .A1(n2389), .A2(n633), .B(n840), .Z(n2392) );
  HDOAI21M20DL U3058 ( .A1(n2189), .A2(n2145), .B(n2025), .Z(n2026) );
  HDOAI21M20DL U3059 ( .A1(n2375), .A2(n2189), .B(n2331), .Z(n2041) );
  HDOAI31DL U3060 ( .A1(n2236), .A2(n2231), .A3(n2211), .B(n2323), .Z(n2150)
         );
  HDAOI21M20DL U3061 ( .A1(n2231), .A2(instruction[26]), .B(n2948), .Z(n2232)
         );
  HDNAN4DL U3062 ( .A1(n2818), .A2(n2817), .A3(n2816), .A4(n2815), .Z(n2823)
         );
  HDAOI21M20DL U3063 ( .A1(n2971), .A2(n2274), .B(n2108), .Z(n2071) );
  HDAOI21M20DL U3064 ( .A1(n2339), .A2(n1687), .B(n2337), .Z(n2369) );
  HDNAN4DL U3065 ( .A1(n2511), .A2(n2254), .A3(n2889), .A4(n2483), .Z(n2206)
         );
  HDNAN3DL U3066 ( .A1(n2851), .A2(n2524), .A3(n2582), .Z(n2172) );
  HDAOI21M20DL U3067 ( .A1(n2212), .A2(n2211), .B(n1704), .Z(n2224) );
  HDNAN3DL U3068 ( .A1(n2778), .A2(n1685), .A3(n1599), .Z(n2779) );
  HDOAI21M20DL U3069 ( .A1(n2107), .A2(n2732), .B(n1686), .Z(n2088) );
  HDOAI222DL U3070 ( .A1(n2244), .A2(n2377), .B1(n2243), .B2(n2033), .C1(n2578), .C2(n2032), .Z(n2036) );
  HDOAI22DL U3071 ( .A1(instruction[25]), .A2(n1704), .B1(n2619), .B2(n2578), 
        .Z(n2153) );
  HDOAI21M20DL U3072 ( .A1(n2668), .A2(n1701), .B(n2694), .Z(n2669) );
  HDOAI21M20DL U3073 ( .A1(n2723), .A2(n1549), .B(n2719), .Z(n1798) );
  HDNAN2D2 U3074 ( .A1(instruction[23]), .A2(instruction[24]), .Z(n1740) );
endmodule

