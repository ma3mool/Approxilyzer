
module sparc_exu_alu ( so, alu_byp_rd_data_e, exu_ifu_brpc_e, 
        exu_lsu_ldst_va_e, exu_lsu_early_va_e, exu_mmu_early_va_e, 
        alu_ecl_add_n64_e, alu_ecl_add_n32_e, alu_ecl_log_n64_e, 
        alu_ecl_log_n32_e, alu_ecl_zhigh_e, alu_ecl_zlow_e, exu_ifu_regz_e, 
        exu_ifu_regn_e, alu_ecl_adderin2_63_e, alu_ecl_adderin2_31_e, 
        alu_ecl_adder_out_63_e, alu_ecl_cout32_e, alu_ecl_cout64_e_l, 
        alu_ecl_mem_addr_invalid_e_l, rclk, se, si, byp_alu_rs1_data_e, 
        byp_alu_rs2_data_e_l, byp_alu_rs3_data_e, byp_alu_rcc_data_e, 
        ecl_alu_cin_e, ifu_exu_invert_d, ecl_alu_log_sel_and_e, 
        ecl_alu_log_sel_or_e, ecl_alu_log_sel_xor_e, ecl_alu_log_sel_move_e, 
        ecl_alu_out_sel_sum_e_l, ecl_alu_out_sel_rs3_e_l, 
        ecl_alu_out_sel_shift_e_l, ecl_alu_out_sel_logic_e_l, 
        shft_alu_shift_out_e, ecl_alu_sethi_inst_e, ifu_lsu_casa_e );
  output [63:0] alu_byp_rd_data_e;
  output [47:0] exu_ifu_brpc_e;
  output [47:0] exu_lsu_ldst_va_e;
  output [10:3] exu_lsu_early_va_e;
  output [7:0] exu_mmu_early_va_e;
  input [63:0] byp_alu_rs1_data_e;
  input [63:0] byp_alu_rs2_data_e_l;
  input [63:0] byp_alu_rs3_data_e;
  input [63:0] byp_alu_rcc_data_e;
  input [63:0] shft_alu_shift_out_e;
  input rclk, se, si, ecl_alu_cin_e, ifu_exu_invert_d, ecl_alu_log_sel_and_e,
         ecl_alu_log_sel_or_e, ecl_alu_log_sel_xor_e, ecl_alu_log_sel_move_e,
         ecl_alu_out_sel_sum_e_l, ecl_alu_out_sel_rs3_e_l,
         ecl_alu_out_sel_shift_e_l, ecl_alu_out_sel_logic_e_l,
         ecl_alu_sethi_inst_e, ifu_lsu_casa_e;
  output so, alu_ecl_add_n64_e, alu_ecl_add_n32_e, alu_ecl_log_n64_e,
         alu_ecl_log_n32_e, alu_ecl_zhigh_e, alu_ecl_zlow_e, exu_ifu_regz_e,
         exu_ifu_regn_e, alu_ecl_adderin2_63_e, alu_ecl_adderin2_31_e,
         alu_ecl_adder_out_63_e, alu_ecl_cout32_e, alu_ecl_cout64_e_l,
         alu_ecl_mem_addr_invalid_e_l;
  wire   exu_ifu_brpc_e_31_, alu_ecl_adder_out_63_e, byp_alu_rcc_data_e_63_,
         invert_e, addsub_cout64_e, addsub_rs2_data_0, addsub_rs2_data_1,
         addsub_rs2_data_2, addsub_rs2_data_3, addsub_rs2_data_4,
         addsub_rs2_data_5, addsub_rs2_data_6, addsub_rs2_data_7,
         addsub_rs2_data_8, addsub_rs2_data_9, addsub_rs2_data_10,
         addsub_rs2_data_11, addsub_rs2_data_12, addsub_rs2_data_13,
         addsub_rs2_data_14, addsub_rs2_data_15, addsub_rs2_data_16,
         addsub_rs2_data_17, addsub_rs2_data_18, addsub_rs2_data_19,
         addsub_rs2_data_20, addsub_rs2_data_21, addsub_rs2_data_22,
         addsub_rs2_data_23, addsub_rs2_data_24, addsub_rs2_data_25,
         addsub_rs2_data_26, addsub_rs2_data_27, addsub_rs2_data_28,
         addsub_rs2_data_29, addsub_rs2_data_30, addsub_rs2_data_32_,
         addsub_rs2_data_33_, addsub_rs2_data_34_, addsub_rs2_data_35_,
         addsub_rs2_data_36_, addsub_rs2_data_37_, addsub_rs2_data_38_,
         addsub_rs2_data_39_, addsub_rs2_data_40_, addsub_rs2_data_41_,
         addsub_rs2_data_42_, addsub_rs2_data_43_, addsub_rs2_data_44_,
         addsub_rs2_data_45_, addsub_rs2_data_46_, addsub_rs2_data_47_,
         addsub_rs2_data_48_, addsub_rs2_data_49_, addsub_rs2_data_50_,
         addsub_rs2_data_51_, addsub_rs2_data_52_, addsub_rs2_data_53_,
         addsub_rs2_data_54_, addsub_rs2_data_55_, addsub_rs2_data_56_,
         addsub_rs2_data_57_, addsub_rs2_data_58_, addsub_rs2_data_59_,
         addsub_rs2_data_60_, addsub_rs2_data_61_, addsub_rs2_data_62_, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n265, n266, n267, n268, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n414, n415, n417, n418, n419, n420, n421, n422, n425, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n873,
         n875, n880, n881, n882, n883, n884, n885, n894, n895, n896, n902,
         n903, n904, n905, n907, n908, n909, n910, n911, n912, n913, n921,
         n923, n927, n928, n929, addsub_adder_add_24_2_DP_OP_276_5026_1_n65,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n64,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n63,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n62,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n61,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n60,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n59,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n58,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n57,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n56,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n55,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n54,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n53,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n52,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n51,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n50,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n49,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n48,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n47,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n46,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n45,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n44,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n43,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n42,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n41,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n40,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n39,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n38,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n37,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n36,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n35,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n32,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n31,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n30,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n29,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n28,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n27,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n26,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n25,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n24,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n23,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n22,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n21,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n20,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n19,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n18,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n17,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n16,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n15,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n14,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n13,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n12,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n11,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n10,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n9,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n8,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n7,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n6,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n5,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n4,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n3,
         addsub_adder_add_24_2_DP_OP_276_5026_1_n2, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968;
  wire   [62:48] adder_out;
  wire   [0:63] addsub_subtract_e;
  assign alu_ecl_add_n32_e = exu_ifu_brpc_e_31_;
  assign exu_ifu_brpc_e[31] = exu_ifu_brpc_e_31_;
  assign exu_ifu_brpc_e[10] = exu_lsu_early_va_e[10];
  assign exu_ifu_brpc_e[9] = exu_lsu_early_va_e[9];
  assign exu_ifu_brpc_e[8] = exu_lsu_early_va_e[8];
  assign exu_mmu_early_va_e[7] = exu_lsu_early_va_e[7];
  assign exu_ifu_brpc_e[7] = exu_lsu_early_va_e[7];
  assign exu_mmu_early_va_e[6] = exu_lsu_early_va_e[6];
  assign exu_ifu_brpc_e[6] = exu_lsu_early_va_e[6];
  assign exu_mmu_early_va_e[5] = exu_lsu_early_va_e[5];
  assign exu_ifu_brpc_e[5] = exu_lsu_early_va_e[5];
  assign exu_mmu_early_va_e[4] = exu_lsu_early_va_e[4];
  assign exu_ifu_brpc_e[4] = exu_lsu_early_va_e[4];
  assign exu_mmu_early_va_e[3] = exu_lsu_early_va_e[3];
  assign exu_ifu_brpc_e[3] = exu_lsu_early_va_e[3];
  assign exu_ifu_brpc_e[2] = exu_mmu_early_va_e[2];
  assign exu_ifu_brpc_e[1] = exu_mmu_early_va_e[1];
  assign exu_ifu_brpc_e[0] = exu_mmu_early_va_e[0];
  assign alu_ecl_add_n64_e = alu_ecl_adder_out_63_e;
  assign exu_ifu_regn_e = byp_alu_rcc_data_e_63_;
  assign byp_alu_rcc_data_e_63_ = byp_alu_rcc_data_e[63];

  HDDFFPQ1 addsub_sub_dff_q_reg_0_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[0]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_1_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[1]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_2_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[2]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_3_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[3]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_4_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[4]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_5_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[5]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_6_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[6]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_7_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[7]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_8_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[8]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_9_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[9]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_10_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[10]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_11_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[11]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_12_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[12]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_13_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[13]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_14_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[14]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_15_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[15]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_16_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[16]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_17_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[17]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_18_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[18]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_19_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[19]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_20_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[20]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_21_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[21]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_22_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[22]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_23_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[23]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_24_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[24]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_25_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[25]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_26_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[26]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_27_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[27]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_28_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[28]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_29_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[29]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_30_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[30]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_31_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[31]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_32_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[32]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_33_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[33]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_34_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[34]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_35_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[35]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_36_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[36]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_37_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[37]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_38_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[38]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_39_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[39]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_40_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[40]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_41_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[41]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_42_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[42]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_43_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[43]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_44_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[44]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_45_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[45]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_46_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[46]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_47_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[47]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_48_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[48]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_49_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[49]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_50_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[50]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_51_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[51]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_52_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[52]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_53_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[53]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_54_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[54]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_55_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[55]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_56_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[56]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_57_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[57]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_58_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[58]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_59_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[59]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_60_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[60]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_61_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[61]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_62_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[62]) );
  HDDFFPQ1 addsub_sub_dff_q_reg_63_ ( .D(n953), .CK(rclk), .Q(
        addsub_subtract_e[63]) );
  HDMUXB2DL U566 ( .A0(byp_alu_rs2_data_e_l[59]), .A1(n902), .SL(
        addsub_subtract_e[59]), .Z(addsub_rs2_data_59_) );
  HDMUXB2DL U568 ( .A0(byp_alu_rs2_data_e_l[58]), .A1(n903), .SL(
        addsub_subtract_e[58]), .Z(addsub_rs2_data_58_) );
  HDMUXB2DL U570 ( .A0(byp_alu_rs2_data_e_l[57]), .A1(n904), .SL(
        addsub_subtract_e[57]), .Z(addsub_rs2_data_57_) );
  HDMUXB2DL U572 ( .A0(byp_alu_rs2_data_e_l[56]), .A1(n905), .SL(
        addsub_subtract_e[56]), .Z(addsub_rs2_data_56_) );
  HDMUXB2DL U576 ( .A0(byp_alu_rs2_data_e_l[54]), .A1(n907), .SL(
        addsub_subtract_e[54]), .Z(addsub_rs2_data_54_) );
  HDMUXB2DL U578 ( .A0(byp_alu_rs2_data_e_l[53]), .A1(n908), .SL(
        addsub_subtract_e[53]), .Z(addsub_rs2_data_53_) );
  HDMUXB2DL U580 ( .A0(byp_alu_rs2_data_e_l[52]), .A1(n909), .SL(
        addsub_subtract_e[52]), .Z(addsub_rs2_data_52_) );
  HDMUXB2DL U582 ( .A0(byp_alu_rs2_data_e_l[51]), .A1(n910), .SL(
        addsub_subtract_e[51]), .Z(addsub_rs2_data_51_) );
  HDMUXB2DL U584 ( .A0(byp_alu_rs2_data_e_l[50]), .A1(n911), .SL(
        addsub_subtract_e[50]), .Z(addsub_rs2_data_50_) );
  HDMUXB2DL U586 ( .A0(byp_alu_rs2_data_e_l[49]), .A1(n912), .SL(
        addsub_subtract_e[49]), .Z(addsub_rs2_data_49_) );
  HDMUXB2DL U588 ( .A0(byp_alu_rs2_data_e_l[48]), .A1(n913), .SL(
        addsub_subtract_e[48]), .Z(addsub_rs2_data_48_) );
  HDMUXB2DL U101 ( .A0(adder_out[60]), .A1(byp_alu_rs1_data_e[60]), .SL(
        ifu_lsu_casa_e), .Z(n382) );
  HDMUXB2DL U100 ( .A0(adder_out[62]), .A1(byp_alu_rs1_data_e[62]), .SL(
        ifu_lsu_casa_e), .Z(n390) );
  HDMUXB2DL U99 ( .A0(n382), .A1(n407), .SL(n390), .Z(n408) );
  HDMUXB2DL U98 ( .A0(adder_out[48]), .A1(byp_alu_rs1_data_e[48]), .SL(
        ifu_lsu_casa_e), .Z(n403) );
  HDMUXB2DL U97 ( .A0(adder_out[59]), .A1(byp_alu_rs1_data_e[59]), .SL(
        ifu_lsu_casa_e), .Z(n383) );
  HDMUXB2DL U96 ( .A0(adder_out[58]), .A1(byp_alu_rs1_data_e[58]), .SL(
        ifu_lsu_casa_e), .Z(n388) );
  HDEXOR2DL U95 ( .A1(n383), .A2(n388), .Z(n410) );
  HDMUXB2DL U93 ( .A0(adder_out[53]), .A1(byp_alu_rs1_data_e[53]), .SL(
        ifu_lsu_casa_e), .Z(n398) );
  HDMUXB2DL U91 ( .A0(adder_out[52]), .A1(byp_alu_rs1_data_e[52]), .SL(
        ifu_lsu_casa_e), .Z(n401) );
  HDMUXB2DL U89 ( .A0(adder_out[51]), .A1(byp_alu_rs1_data_e[51]), .SL(
        ifu_lsu_casa_e), .Z(n402) );
  HDEXOR2DL U88 ( .A1(n402), .A2(n393), .Z(n406) );
  HDMUXB2DL U87 ( .A0(adder_out[49]), .A1(byp_alu_rs1_data_e[49]), .SL(
        ifu_lsu_casa_e), .Z(n392) );
  HDMUXB2DL U86 ( .A0(n392), .A1(n393), .SL(n403), .Z(n394) );
  HDMUXB2DL U85 ( .A0(adder_out[56]), .A1(byp_alu_rs1_data_e[56]), .SL(
        ifu_lsu_casa_e), .Z(n386) );
  HDEXNOR2DL U83 ( .A1(n401), .A2(n402), .Z(n400) );
  HDMUXB2DL U81 ( .A0(alu_ecl_adder_out_63_e), .A1(byp_alu_rs1_data_e[63]), 
        .SL(ifu_lsu_casa_e), .Z(n391) );
  HDEXNOR2DL U80 ( .A1(n390), .A2(n391), .Z(n378) );
  HDMUXB2DL U79 ( .A0(adder_out[57]), .A1(byp_alu_rs1_data_e[57]), .SL(
        ifu_lsu_casa_e), .Z(n387) );
  HDEXNOR2DL U77 ( .A1(n384), .A2(n385), .Z(n380) );
  HDEXNOR2DL U76 ( .A1(n382), .A2(n383), .Z(n381) );
  HDMUXB2DL U430 ( .A0(invert_e), .A1(n955), .SL(byp_alu_rs2_data_e_l[19]), 
        .Z(n796) );
  HDAO32DL U426 ( .A1(n796), .A2(n127), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n796), .Z(n795) );
  HDMUXB2DL U418 ( .A0(invert_e), .A1(n956), .SL(byp_alu_rs2_data_e_l[20]), 
        .Z(n782) );
  HDAO32DL U414 ( .A1(n782), .A2(n129), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n782), .Z(n781) );
  HDMUXB2DL U412 ( .A0(invert_e), .A1(n7), .SL(byp_alu_rs2_data_e_l[21]), .Z(
        n775) );
  HDAO32DL U408 ( .A1(n775), .A2(n126), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n775), .Z(n774) );
  HDMUXB2DL U406 ( .A0(n954), .A1(n955), .SL(byp_alu_rs2_data_e_l[22]), .Z(
        n768) );
  HDAO32DL U402 ( .A1(n768), .A2(n136), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n768), .Z(n767) );
  HDMUXB2DL U454 ( .A0(n954), .A1(n956), .SL(byp_alu_rs2_data_e_l[15]), .Z(
        n824) );
  HDAO32DL U450 ( .A1(n824), .A2(n121), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n824), .Z(n823) );
  HDMUXB2DL U448 ( .A0(n954), .A1(n955), .SL(byp_alu_rs2_data_e_l[16]), .Z(
        n817) );
  HDAO32DL U444 ( .A1(n817), .A2(n119), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n817), .Z(n816) );
  HDMUXB2DL U442 ( .A0(n954), .A1(n7), .SL(byp_alu_rs2_data_e_l[17]), .Z(n810)
         );
  HDAO32DL U438 ( .A1(n810), .A2(n120), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n810), .Z(n809) );
  HDMUXB2DL U436 ( .A0(invert_e), .A1(n956), .SL(byp_alu_rs2_data_e_l[18]), 
        .Z(n803) );
  HDAO32DL U432 ( .A1(n803), .A2(n128), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n803), .Z(n802) );
  HDMUXB2DL U376 ( .A0(invert_e), .A1(n956), .SL(byp_alu_rs2_data_e_l[27]), 
        .Z(n733) );
  HDAO32DL U372 ( .A1(n733), .A2(n147), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n733), .Z(n732) );
  HDMUXB2DL U370 ( .A0(invert_e), .A1(n955), .SL(byp_alu_rs2_data_e_l[28]), 
        .Z(n726) );
  HDAO32DL U366 ( .A1(n726), .A2(n145), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n726), .Z(n725) );
  HDMUXB2DL U364 ( .A0(invert_e), .A1(n7), .SL(byp_alu_rs2_data_e_l[29]), .Z(
        n719) );
  HDAO32DL U360 ( .A1(n719), .A2(n146), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n719), .Z(n718) );
  HDMUXB2DL U352 ( .A0(invert_e), .A1(n956), .SL(byp_alu_rs2_data_e_l[30]), 
        .Z(n705) );
  HDAO32DL U348 ( .A1(n705), .A2(n148), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n705), .Z(n704) );
  HDMUXB2DL U400 ( .A0(invert_e), .A1(n7), .SL(byp_alu_rs2_data_e_l[23]), .Z(
        n761) );
  HDAO32DL U396 ( .A1(n761), .A2(n135), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n761), .Z(n760) );
  HDMUXB2DL U394 ( .A0(invert_e), .A1(n955), .SL(byp_alu_rs2_data_e_l[24]), 
        .Z(n754) );
  HDAO32DL U390 ( .A1(n754), .A2(n137), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n754), .Z(n753) );
  HDMUXB2DL U388 ( .A0(invert_e), .A1(n7), .SL(byp_alu_rs2_data_e_l[25]), .Z(
        n747) );
  HDAO32DL U384 ( .A1(n747), .A2(n138), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n747), .Z(n746) );
  HDMUXB2DL U382 ( .A0(invert_e), .A1(n955), .SL(byp_alu_rs2_data_e_l[26]), 
        .Z(n740) );
  HDAO32DL U378 ( .A1(n740), .A2(n134), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n740), .Z(n739) );
  HDMUXB2DL U292 ( .A0(invert_e), .A1(n955), .SL(byp_alu_rs2_data_e_l[3]), .Z(
        n635) );
  HDAO32DL U288 ( .A1(n635), .A2(n85), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n635), .Z(n634) );
  HDMUXB2DL U226 ( .A0(invert_e), .A1(n955), .SL(byp_alu_rs2_data_e_l[4]), .Z(
        n558) );
  HDAO32DL U222 ( .A1(n558), .A2(n160), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n558), .Z(n557) );
  HDMUXB2DL U160 ( .A0(invert_e), .A1(n956), .SL(byp_alu_rs2_data_e_l[5]), .Z(
        n481) );
  HDAO32DL U156 ( .A1(n481), .A2(n157), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n481), .Z(n480) );
  HDMUXB2DL U130 ( .A0(invert_e), .A1(n7), .SL(byp_alu_rs2_data_e_l[6]), .Z(
        n446) );
  HDAO32DL U126 ( .A1(n446), .A2(n159), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n446), .Z(n445) );
  HDMUXB2DL U346 ( .A0(invert_e), .A1(n7), .SL(byp_alu_rs2_data_e_l[31]), .Z(
        n698) );
  HDMUXB2DL U495 ( .A0(n954), .A1(n7), .SL(byp_alu_rs2_data_e_l[0]), .Z(n866)
         );
  HDAO32DL U489 ( .A1(n866), .A2(n86), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n866), .Z(n865) );
  HDMUXB2DL U424 ( .A0(invert_e), .A1(n956), .SL(byp_alu_rs2_data_e_l[1]), .Z(
        n789) );
  HDAO32DL U420 ( .A1(n789), .A2(n80), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n789), .Z(n788) );
  HDMUXB2DL U358 ( .A0(invert_e), .A1(n955), .SL(byp_alu_rs2_data_e_l[2]), .Z(
        n712) );
  HDAO32DL U354 ( .A1(n712), .A2(n81), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n712), .Z(n711) );
  HDMUXB2DL U478 ( .A0(n954), .A1(n7), .SL(byp_alu_rs2_data_e_l[11]), .Z(n852)
         );
  HDAO32DL U474 ( .A1(n852), .A2(n110), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n852), .Z(n851) );
  HDMUXB2DL U472 ( .A0(n954), .A1(n7), .SL(byp_alu_rs2_data_e_l[12]), .Z(n845)
         );
  HDAO32DL U468 ( .A1(n845), .A2(n153), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n845), .Z(n844) );
  HDMUXB2DL U466 ( .A0(n954), .A1(n7), .SL(byp_alu_rs2_data_e_l[13]), .Z(n838)
         );
  HDAO32DL U462 ( .A1(n838), .A2(n107), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n838), .Z(n837) );
  HDMUXB2DL U460 ( .A0(n954), .A1(n955), .SL(byp_alu_rs2_data_e_l[14]), .Z(
        n831) );
  HDAO32DL U456 ( .A1(n831), .A2(n108), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n831), .Z(n830) );
  HDMUXB2DL U124 ( .A0(invert_e), .A1(n7), .SL(byp_alu_rs2_data_e_l[7]), .Z(
        n439) );
  HDAO32DL U120 ( .A1(n439), .A2(n155), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n439), .Z(n438) );
  HDMUXB2DL U118 ( .A0(invert_e), .A1(n7), .SL(byp_alu_rs2_data_e_l[8]), .Z(
        n432) );
  HDAO32DL U114 ( .A1(n432), .A2(n156), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n432), .Z(n431) );
  HDMUXB2DL U112 ( .A0(invert_e), .A1(n7), .SL(byp_alu_rs2_data_e_l[9]), .Z(
        n421) );
  HDAO32DL U108 ( .A1(n421), .A2(n158), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n421), .Z(n420) );
  HDMUXB2DL U484 ( .A0(n954), .A1(n7), .SL(byp_alu_rs2_data_e_l[10]), .Z(n859)
         );
  HDAO32DL U480 ( .A1(n859), .A2(n154), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n859), .Z(n858) );
  HDMUXB2DL U39 ( .A0(byp_alu_rs1_data_e[4]), .A1(n160), .SL(addsub_rs2_data_4), .Z(n51) );
  HDMUXB2DL U38 ( .A0(byp_alu_rs1_data_e[6]), .A1(n159), .SL(addsub_rs2_data_6), .Z(n43) );
  HDMUXB2DL U37 ( .A0(byp_alu_rs1_data_e[9]), .A1(n158), .SL(addsub_rs2_data_9), .Z(n39) );
  HDMUXB2DL U36 ( .A0(byp_alu_rs1_data_e[5]), .A1(n157), .SL(addsub_rs2_data_5), .Z(n49) );
  HDMUXB2DL U35 ( .A0(byp_alu_rs1_data_e[8]), .A1(n156), .SL(addsub_rs2_data_8), .Z(n42) );
  HDMUXB2DL U34 ( .A0(byp_alu_rs1_data_e[7]), .A1(n155), .SL(addsub_rs2_data_7), .Z(n44) );
  HDMUXB2DL U33 ( .A0(byp_alu_rs1_data_e[10]), .A1(n154), .SL(
        addsub_rs2_data_10), .Z(n41) );
  HDMUXB2DL U32 ( .A0(byp_alu_rs1_data_e[12]), .A1(n153), .SL(
        addsub_rs2_data_12), .Z(n70) );
  HDMUXB2DL U31 ( .A0(byp_alu_rs1_data_e[30]), .A1(n148), .SL(
        addsub_rs2_data_30), .Z(n63) );
  HDMUXB2DL U30 ( .A0(byp_alu_rs1_data_e[27]), .A1(n147), .SL(
        addsub_rs2_data_27), .Z(n93) );
  HDMUXB2DL U29 ( .A0(byp_alu_rs1_data_e[29]), .A1(n146), .SL(
        addsub_rs2_data_29), .Z(n61) );
  HDMUXB2DL U28 ( .A0(byp_alu_rs1_data_e[28]), .A1(n145), .SL(
        addsub_rs2_data_28), .Z(n62) );
  HDMUXB2DL U27 ( .A0(n143), .A1(byp_alu_rs1_data_e[31]), .SL(n144), .Z(n60)
         );
  HDMUXB2DL U26 ( .A0(byp_alu_rs1_data_e[25]), .A1(n138), .SL(
        addsub_rs2_data_25), .Z(n92) );
  HDMUXB2DL U25 ( .A0(byp_alu_rs1_data_e[24]), .A1(n137), .SL(
        addsub_rs2_data_24), .Z(n96) );
  HDMUXB2DL U24 ( .A0(byp_alu_rs1_data_e[22]), .A1(n136), .SL(
        addsub_rs2_data_22), .Z(n95) );
  HDMUXB2DL U23 ( .A0(byp_alu_rs1_data_e[23]), .A1(n135), .SL(
        addsub_rs2_data_23), .Z(n94) );
  HDMUXB2DL U22 ( .A0(byp_alu_rs1_data_e[26]), .A1(n134), .SL(
        addsub_rs2_data_26), .Z(n91) );
  HDMUXB2DL U21 ( .A0(byp_alu_rs1_data_e[20]), .A1(n129), .SL(
        addsub_rs2_data_20), .Z(n97) );
  HDMUXB2DL U20 ( .A0(byp_alu_rs1_data_e[18]), .A1(n128), .SL(
        addsub_rs2_data_18), .Z(n106) );
  HDMUXB2DL U19 ( .A0(byp_alu_rs1_data_e[19]), .A1(n127), .SL(
        addsub_rs2_data_19), .Z(n98) );
  HDMUXB2DL U18 ( .A0(byp_alu_rs1_data_e[21]), .A1(n126), .SL(
        addsub_rs2_data_21), .Z(n103) );
  HDMUXB2DL U17 ( .A0(byp_alu_rs1_data_e[15]), .A1(n121), .SL(
        addsub_rs2_data_15), .Z(n109) );
  HDMUXB2DL U16 ( .A0(byp_alu_rs1_data_e[17]), .A1(n120), .SL(
        addsub_rs2_data_17), .Z(n104) );
  HDMUXB2DL U15 ( .A0(byp_alu_rs1_data_e[16]), .A1(n119), .SL(
        addsub_rs2_data_16), .Z(n105) );
  HDMUXB2DL U14 ( .A0(byp_alu_rs1_data_e[11]), .A1(n110), .SL(
        addsub_rs2_data_11), .Z(n40) );
  HDMUXB2DL U13 ( .A0(byp_alu_rs1_data_e[14]), .A1(n108), .SL(
        addsub_rs2_data_14), .Z(n69) );
  HDMUXB2DL U12 ( .A0(byp_alu_rs1_data_e[13]), .A1(n107), .SL(
        addsub_rs2_data_13), .Z(n68) );
  HDMUXB2DL U11 ( .A0(byp_alu_rs1_data_e[0]), .A1(n86), .SL(ecl_alu_cin_e), 
        .Z(n82) );
  HDMUXB2DL U9 ( .A0(byp_alu_rs1_data_e[3]), .A1(n85), .SL(addsub_rs2_data_3), 
        .Z(n50) );
  HDMUXB2DL U8 ( .A0(byp_alu_rs1_data_e[2]), .A1(n81), .SL(addsub_rs2_data_2), 
        .Z(n52) );
  HDMUXB2DL U7 ( .A0(byp_alu_rs1_data_e[1]), .A1(n80), .SL(addsub_rs2_data_1), 
        .Z(n71) );
  HDMUXB2DL U214 ( .A0(invert_e), .A1(n7), .SL(byp_alu_rs2_data_e_l[51]), .Z(
        n544) );
  HDAO32DL U210 ( .A1(n544), .A2(n282), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n544), .Z(n543) );
  HDMUXB2DL U208 ( .A0(invert_e), .A1(n7), .SL(byp_alu_rs2_data_e_l[52]), .Z(
        n537) );
  HDAO32DL U204 ( .A1(n537), .A2(n284), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n537), .Z(n536) );
  HDMUXB2DL U202 ( .A0(invert_e), .A1(n956), .SL(byp_alu_rs2_data_e_l[53]), 
        .Z(n530) );
  HDAO32DL U198 ( .A1(n530), .A2(n280), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n530), .Z(n529) );
  HDMUXB2DL U196 ( .A0(invert_e), .A1(n955), .SL(byp_alu_rs2_data_e_l[54]), 
        .Z(n523) );
  HDAO32DL U192 ( .A1(n523), .A2(n281), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n523), .Z(n522) );
  HDMUXB2DL U244 ( .A0(invert_e), .A1(n956), .SL(byp_alu_rs2_data_e_l[47]), 
        .Z(n579) );
  HDAO32DL U240 ( .A1(n579), .A2(n311), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n579), .Z(n578) );
  HDMUXB2DL U238 ( .A0(invert_e), .A1(n7), .SL(byp_alu_rs2_data_e_l[48]), .Z(
        n572) );
  HDAO32DL U234 ( .A1(n572), .A2(n309), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n572), .Z(n571) );
  HDMUXB2DL U232 ( .A0(invert_e), .A1(n7), .SL(byp_alu_rs2_data_e_l[49]), .Z(
        n565) );
  HDAO32DL U228 ( .A1(n565), .A2(n291), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n565), .Z(n564) );
  HDMUXB2DL U220 ( .A0(invert_e), .A1(n955), .SL(byp_alu_rs2_data_e_l[50]), 
        .Z(n551) );
  HDAO32DL U216 ( .A1(n551), .A2(n285), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n551), .Z(n550) );
  HDMUXB2DL U166 ( .A0(invert_e), .A1(n955), .SL(byp_alu_rs2_data_e_l[59]), 
        .Z(n488) );
  HDAO32DL U162 ( .A1(n488), .A2(n265), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n488), .Z(n487) );
  HDMUXB2DL U154 ( .A0(invert_e), .A1(n7), .SL(byp_alu_rs2_data_e_l[60]), .Z(
        n474) );
  HDAO32DL U150 ( .A1(n474), .A2(n266), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n474), .Z(n473) );
  HDMUXB2DL U148 ( .A0(invert_e), .A1(n955), .SL(byp_alu_rs2_data_e_l[61]), 
        .Z(n467) );
  HDAO32DL U144 ( .A1(n467), .A2(n268), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n467), .Z(n466) );
  HDMUXB2DL U142 ( .A0(invert_e), .A1(n956), .SL(byp_alu_rs2_data_e_l[62]), 
        .Z(n460) );
  HDAO32DL U138 ( .A1(n460), .A2(n270), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n460), .Z(n459) );
  HDMUXB2DL U190 ( .A0(invert_e), .A1(n7), .SL(byp_alu_rs2_data_e_l[55]), .Z(
        n516) );
  HDAO32DL U186 ( .A1(n516), .A2(n283), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n516), .Z(n515) );
  HDMUXB2DL U184 ( .A0(invert_e), .A1(n7), .SL(byp_alu_rs2_data_e_l[56]), .Z(
        n509) );
  HDAO32DL U180 ( .A1(n509), .A2(n275), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n509), .Z(n508) );
  HDMUXB2DL U178 ( .A0(invert_e), .A1(n956), .SL(byp_alu_rs2_data_e_l[57]), 
        .Z(n502) );
  HDAO32DL U174 ( .A1(n502), .A2(n267), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n502), .Z(n501) );
  HDMUXB2DL U172 ( .A0(invert_e), .A1(n7), .SL(byp_alu_rs2_data_e_l[58]), .Z(
        n495) );
  HDAO32DL U168 ( .A1(n495), .A2(n271), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n495), .Z(n494) );
  HDMUXB2DL U322 ( .A0(invert_e), .A1(n7), .SL(byp_alu_rs2_data_e_l[35]), .Z(
        n670) );
  HDAO32DL U318 ( .A1(n670), .A2(n333), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n670), .Z(n669) );
  HDMUXB2DL U316 ( .A0(invert_e), .A1(n7), .SL(byp_alu_rs2_data_e_l[36]), .Z(
        n663) );
  HDAO32DL U312 ( .A1(n663), .A2(n332), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n663), .Z(n662) );
  HDMUXB2DL U310 ( .A0(invert_e), .A1(n956), .SL(byp_alu_rs2_data_e_l[37]), 
        .Z(n656) );
  HDAO32DL U306 ( .A1(n656), .A2(n331), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n656), .Z(n655) );
  HDMUXB2DL U304 ( .A0(invert_e), .A1(n955), .SL(byp_alu_rs2_data_e_l[38]), 
        .Z(n649) );
  HDAO32DL U300 ( .A1(n649), .A2(n330), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n649), .Z(n648) );
  HDMUXB2DL U136 ( .A0(invert_e), .A1(n956), .SL(byp_alu_rs2_data_e_l[63]), 
        .Z(n453) );
  HDMUXB2DL U135 ( .A0(ecl_alu_log_sel_xor_e), .A1(ecl_alu_log_sel_and_e), 
        .SL(n453), .Z(n454) );
  HDOAI21M20DL U134 ( .A1(n968), .A2(n454), .B(byp_alu_rs1_data_e[63]), .Z(
        n451) );
  HDMUXB2DL U340 ( .A0(invert_e), .A1(n956), .SL(byp_alu_rs2_data_e_l[32]), 
        .Z(n691) );
  HDAO32DL U336 ( .A1(n691), .A2(n315), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n691), .Z(n690) );
  HDMUXB2DL U334 ( .A0(invert_e), .A1(n956), .SL(byp_alu_rs2_data_e_l[33]), 
        .Z(n684) );
  HDAO32DL U330 ( .A1(n684), .A2(n314), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n684), .Z(n683) );
  HDMUXB2DL U328 ( .A0(n954), .A1(n955), .SL(byp_alu_rs2_data_e_l[34]), .Z(
        n677) );
  HDAO32DL U324 ( .A1(n677), .A2(n313), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n677), .Z(n676) );
  HDMUXB2DL U268 ( .A0(invert_e), .A1(n956), .SL(byp_alu_rs2_data_e_l[43]), 
        .Z(n607) );
  HDAO32DL U264 ( .A1(n607), .A2(n321), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n607), .Z(n606) );
  HDMUXB2DL U262 ( .A0(invert_e), .A1(n7), .SL(byp_alu_rs2_data_e_l[44]), .Z(
        n600) );
  HDAO32DL U258 ( .A1(n600), .A2(n320), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n600), .Z(n599) );
  HDMUXB2DL U256 ( .A0(invert_e), .A1(n7), .SL(byp_alu_rs2_data_e_l[45]), .Z(
        n593) );
  HDAO32DL U252 ( .A1(n593), .A2(n312), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n593), .Z(n592) );
  HDMUXB2DL U250 ( .A0(invert_e), .A1(n955), .SL(byp_alu_rs2_data_e_l[46]), 
        .Z(n586) );
  HDAO32DL U246 ( .A1(n586), .A2(n310), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n586), .Z(n585) );
  HDMUXB2DL U298 ( .A0(n954), .A1(n956), .SL(byp_alu_rs2_data_e_l[39]), .Z(
        n642) );
  HDAO32DL U294 ( .A1(n642), .A2(n329), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n642), .Z(n641) );
  HDMUXB2DL U286 ( .A0(invert_e), .A1(n7), .SL(byp_alu_rs2_data_e_l[40]), .Z(
        n628) );
  HDAO32DL U282 ( .A1(n628), .A2(n324), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n628), .Z(n627) );
  HDMUXB2DL U280 ( .A0(invert_e), .A1(n955), .SL(byp_alu_rs2_data_e_l[41]), 
        .Z(n621) );
  HDAO32DL U276 ( .A1(n621), .A2(n323), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n621), .Z(n620) );
  HDMUXB2DL U274 ( .A0(invert_e), .A1(n956), .SL(byp_alu_rs2_data_e_l[42]), 
        .Z(n614) );
  HDAO32DL U270 ( .A1(n614), .A2(n322), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n614), .Z(n613) );
  HDMUXB2DL U75 ( .A0(byp_alu_rs1_data_e[35]), .A1(n333), .SL(
        addsub_rs2_data_35_), .Z(n219) );
  HDMUXB2DL U74 ( .A0(byp_alu_rs1_data_e[36]), .A1(n332), .SL(
        addsub_rs2_data_36_), .Z(n218) );
  HDMUXB2DL U73 ( .A0(byp_alu_rs1_data_e[37]), .A1(n331), .SL(
        addsub_rs2_data_37_), .Z(n220) );
  HDMUXB2DL U72 ( .A0(byp_alu_rs1_data_e[38]), .A1(n330), .SL(
        addsub_rs2_data_38_), .Z(n216) );
  HDMUXB2DL U71 ( .A0(byp_alu_rs1_data_e[39]), .A1(n329), .SL(
        addsub_rs2_data_39_), .Z(n297) );
  HDMUXB2DL U70 ( .A0(byp_alu_rs1_data_e[40]), .A1(n324), .SL(
        addsub_rs2_data_40_), .Z(n217) );
  HDMUXB2DL U69 ( .A0(byp_alu_rs1_data_e[41]), .A1(n323), .SL(
        addsub_rs2_data_41_), .Z(n295) );
  HDMUXB2DL U68 ( .A0(byp_alu_rs1_data_e[42]), .A1(n322), .SL(
        addsub_rs2_data_42_), .Z(n294) );
  HDMUXB2DL U67 ( .A0(byp_alu_rs1_data_e[43]), .A1(n321), .SL(
        addsub_rs2_data_43_), .Z(n296) );
  HDMUXB2DL U66 ( .A0(byp_alu_rs1_data_e[44]), .A1(n320), .SL(
        addsub_rs2_data_44_), .Z(n292) );
  HDMUXB2DL U65 ( .A0(byp_alu_rs1_data_e[32]), .A1(n315), .SL(
        addsub_rs2_data_32_), .Z(n222) );
  HDMUXB2DL U64 ( .A0(byp_alu_rs1_data_e[33]), .A1(n314), .SL(
        addsub_rs2_data_33_), .Z(n221) );
  HDMUXB2DL U63 ( .A0(byp_alu_rs1_data_e[34]), .A1(n313), .SL(
        addsub_rs2_data_34_), .Z(n223) );
  HDMUXB2DL U62 ( .A0(byp_alu_rs1_data_e[45]), .A1(n312), .SL(
        addsub_rs2_data_45_), .Z(n290) );
  HDMUXB2DL U61 ( .A0(byp_alu_rs1_data_e[47]), .A1(n311), .SL(
        addsub_rs2_data_47_), .Z(n252) );
  HDMUXB2DL U60 ( .A0(byp_alu_rs1_data_e[46]), .A1(n310), .SL(
        addsub_rs2_data_46_), .Z(n293) );
  HDMUXB2DL U59 ( .A0(byp_alu_rs1_data_e[48]), .A1(n309), .SL(
        addsub_rs2_data_48_), .Z(n253) );
  HDMUXB2DL U58 ( .A0(byp_alu_rs1_data_e[63]), .A1(n304), .SL(
        alu_ecl_adderin2_63_e), .Z(n244) );
  HDMUXB2DL U56 ( .A0(byp_alu_rs1_data_e[49]), .A1(n291), .SL(
        addsub_rs2_data_49_), .Z(n249) );
  HDMUXB2DL U55 ( .A0(byp_alu_rs1_data_e[50]), .A1(n285), .SL(
        addsub_rs2_data_50_), .Z(n250) );
  HDMUXB2DL U54 ( .A0(byp_alu_rs1_data_e[52]), .A1(n284), .SL(
        addsub_rs2_data_52_), .Z(n260) );
  HDMUXB2DL U53 ( .A0(byp_alu_rs1_data_e[55]), .A1(n283), .SL(
        addsub_rs2_data_55_), .Z(n235) );
  HDMUXB2DL U52 ( .A0(byp_alu_rs1_data_e[51]), .A1(n282), .SL(
        addsub_rs2_data_51_), .Z(n251) );
  HDMUXB2DL U51 ( .A0(byp_alu_rs1_data_e[54]), .A1(n281), .SL(
        addsub_rs2_data_54_), .Z(n259) );
  HDMUXB2DL U50 ( .A0(byp_alu_rs1_data_e[53]), .A1(n280), .SL(
        addsub_rs2_data_53_), .Z(n258) );
  HDMUXB2DL U49 ( .A0(byp_alu_rs1_data_e[56]), .A1(n275), .SL(
        addsub_rs2_data_56_), .Z(n236) );
  HDMUXB2DL U48 ( .A0(byp_alu_rs1_data_e[58]), .A1(n271), .SL(
        addsub_rs2_data_58_), .Z(n234) );
  HDMUXB2DL U45 ( .A0(byp_alu_rs1_data_e[62]), .A1(n270), .SL(
        addsub_rs2_data_62_), .Z(n243) );
  HDMUXB2DL U44 ( .A0(byp_alu_rs1_data_e[61]), .A1(n268), .SL(
        addsub_rs2_data_61_), .Z(n242) );
  HDMUXB2DL U43 ( .A0(byp_alu_rs1_data_e[57]), .A1(n267), .SL(
        addsub_rs2_data_57_), .Z(n237) );
  HDMUXB2DL U42 ( .A0(byp_alu_rs1_data_e[60]), .A1(n266), .SL(
        addsub_rs2_data_60_), .Z(n232) );
  HDMUXB2DL U41 ( .A0(byp_alu_rs1_data_e[59]), .A1(n265), .SL(
        addsub_rs2_data_59_), .Z(n233) );
  HDINVD1 U567 ( .A(byp_alu_rs2_data_e_l[59]), .Z(n902) );
  HDINVD1 U569 ( .A(byp_alu_rs2_data_e_l[58]), .Z(n903) );
  HDINVD1 U571 ( .A(byp_alu_rs2_data_e_l[57]), .Z(n904) );
  HDINVD1 U573 ( .A(byp_alu_rs2_data_e_l[56]), .Z(n905) );
  HDINVD1 U577 ( .A(byp_alu_rs2_data_e_l[54]), .Z(n907) );
  HDINVD1 U579 ( .A(byp_alu_rs2_data_e_l[53]), .Z(n908) );
  HDINVD1 U581 ( .A(byp_alu_rs2_data_e_l[52]), .Z(n909) );
  HDINVD1 U583 ( .A(byp_alu_rs2_data_e_l[51]), .Z(n910) );
  HDINVD1 U585 ( .A(byp_alu_rs2_data_e_l[50]), .Z(n911) );
  HDINVD1 U587 ( .A(byp_alu_rs2_data_e_l[49]), .Z(n912) );
  HDINVD1 U589 ( .A(byp_alu_rs2_data_e_l[48]), .Z(n913) );
  HDINVD1 U605 ( .A(byp_alu_rs2_data_e_l[40]), .Z(n921) );
  HDINVD1 U609 ( .A(byp_alu_rs2_data_e_l[38]), .Z(n923) );
  HDINVD1 U617 ( .A(byp_alu_rs2_data_e_l[34]), .Z(n927) );
  HDINVD1 U619 ( .A(byp_alu_rs2_data_e_l[33]), .Z(n928) );
  HDINVD1 U621 ( .A(byp_alu_rs2_data_e_l[32]), .Z(n929) );
  HDINVD1 U523 ( .A(byp_alu_rs2_data_e_l[25]), .Z(n880) );
  HDINVD1 U525 ( .A(byp_alu_rs2_data_e_l[24]), .Z(n881) );
  HDINVD1 U527 ( .A(byp_alu_rs2_data_e_l[23]), .Z(n882) );
  HDINVD1 U529 ( .A(byp_alu_rs2_data_e_l[22]), .Z(n883) );
  HDINVD1 U531 ( .A(byp_alu_rs2_data_e_l[21]), .Z(n884) );
  HDINVD1 U533 ( .A(byp_alu_rs2_data_e_l[20]), .Z(n885) );
  HDINVD1 U551 ( .A(byp_alu_rs2_data_e_l[12]), .Z(n894) );
  HDINVD1 U553 ( .A(byp_alu_rs2_data_e_l[11]), .Z(n895) );
  HDINVD1 U555 ( .A(byp_alu_rs2_data_e_l[10]), .Z(n896) );
  HDINVD1 U509 ( .A(byp_alu_rs2_data_e_l[4]), .Z(n873) );
  HDINVD1 U513 ( .A(byp_alu_rs2_data_e_l[3]), .Z(n875) );
  HDMUX2D1 U849 ( .A0(adder_out[61]), .A1(byp_alu_rs1_data_e[61]), .SL(
        ifu_lsu_casa_e), .Z(n407) );
  HDMUX2D1 U848 ( .A0(exu_ifu_brpc_e[47]), .A1(byp_alu_rs1_data_e[47]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[47]) );
  HDOAI211D1 U846 ( .A1(n382), .A2(n407), .B(n408), .C(n409), .Z(n374) );
  HDINVD1 U92 ( .A(n398), .Z(n404) );
  HDNAN2D1 U90 ( .A1(n404), .A2(n401), .Z(n405) );
  HDMUX2D1 U845 ( .A0(adder_out[50]), .A1(byp_alu_rs1_data_e[50]), .SL(
        ifu_lsu_casa_e), .Z(n393) );
  HDOAI211D1 U844 ( .A1(n404), .A2(n401), .B(n405), .C(n406), .Z(n375) );
  HDMUX2D1 U843 ( .A0(adder_out[55]), .A1(byp_alu_rs1_data_e[55]), .SL(
        ifu_lsu_casa_e), .Z(n385) );
  HDMUX2D1 U842 ( .A0(adder_out[54]), .A1(byp_alu_rs1_data_e[54]), .SL(
        ifu_lsu_casa_e), .Z(n384) );
  HDNAN2D1 U84 ( .A1(n384), .A2(n398), .Z(n399) );
  HDOAI211D1 U841 ( .A1(n384), .A2(n398), .B(n399), .C(n400), .Z(n396) );
  HDNOR2D1 U82 ( .A1(n386), .A2(n385), .Z(n397) );
  HDAOI211D1 U840 ( .A1(n386), .A2(n385), .B(n396), .C(n397), .Z(n395) );
  HDOAI211D1 U839 ( .A1(n392), .A2(n393), .B(n394), .C(n395), .Z(n376) );
  HDNAN3D1 U78 ( .A1(n388), .A2(n386), .A3(n387), .Z(n389) );
  HDOAI31D1 U838 ( .A1(n386), .A2(n387), .A3(n388), .B(n389), .Z(n379) );
  HDNAN4D1 U837 ( .A1(n378), .A2(n379), .A3(n380), .A4(n381), .Z(n377) );
  HDNOR4D1 U836 ( .A1(n374), .A2(n375), .A3(n376), .A4(n377), .Z(
        alu_ecl_mem_addr_invalid_e_l) );
  HDINVD1 U102 ( .A(addsub_cout64_e), .Z(alu_ecl_cout64_e_l) );
  HDNOR4D1 U689 ( .A1(byp_alu_rcc_data_e[9]), .A2(byp_alu_rcc_data_e[8]), .A3(
        byp_alu_rcc_data_e[7]), .A4(byp_alu_rcc_data_e[6]), .Z(n24) );
  HDNOR4D1 U688 ( .A1(byp_alu_rcc_data_e_63_), .A2(byp_alu_rcc_data_e[62]), 
        .A3(byp_alu_rcc_data_e[61]), .A4(byp_alu_rcc_data_e[60]), .Z(n25) );
  HDNOR4D1 U687 ( .A1(byp_alu_rcc_data_e[5]), .A2(byp_alu_rcc_data_e[59]), 
        .A3(byp_alu_rcc_data_e[58]), .A4(byp_alu_rcc_data_e[57]), .Z(n26) );
  HDNOR4D1 U686 ( .A1(byp_alu_rcc_data_e[56]), .A2(byp_alu_rcc_data_e[55]), 
        .A3(byp_alu_rcc_data_e[54]), .A4(byp_alu_rcc_data_e[53]), .Z(n27) );
  HDNAN4D1 U685 ( .A1(n24), .A2(n25), .A3(n26), .A4(n27), .Z(n8) );
  HDNOR4D1 U684 ( .A1(byp_alu_rcc_data_e[52]), .A2(byp_alu_rcc_data_e[51]), 
        .A3(byp_alu_rcc_data_e[50]), .A4(byp_alu_rcc_data_e[4]), .Z(n20) );
  HDNOR4D1 U683 ( .A1(byp_alu_rcc_data_e[49]), .A2(byp_alu_rcc_data_e[48]), 
        .A3(byp_alu_rcc_data_e[47]), .A4(byp_alu_rcc_data_e[46]), .Z(n21) );
  HDNOR4D1 U682 ( .A1(byp_alu_rcc_data_e[45]), .A2(byp_alu_rcc_data_e[44]), 
        .A3(byp_alu_rcc_data_e[43]), .A4(byp_alu_rcc_data_e[42]), .Z(n22) );
  HDNOR4D1 U681 ( .A1(byp_alu_rcc_data_e[41]), .A2(byp_alu_rcc_data_e[40]), 
        .A3(byp_alu_rcc_data_e[3]), .A4(byp_alu_rcc_data_e[39]), .Z(n23) );
  HDNAN4D1 U680 ( .A1(n20), .A2(n21), .A3(n22), .A4(n23), .Z(n9) );
  HDNOR4D1 U679 ( .A1(byp_alu_rcc_data_e[38]), .A2(byp_alu_rcc_data_e[37]), 
        .A3(byp_alu_rcc_data_e[36]), .A4(byp_alu_rcc_data_e[35]), .Z(n16) );
  HDNOR4D1 U678 ( .A1(byp_alu_rcc_data_e[34]), .A2(byp_alu_rcc_data_e[33]), 
        .A3(byp_alu_rcc_data_e[32]), .A4(byp_alu_rcc_data_e[31]), .Z(n17) );
  HDNOR4D1 U677 ( .A1(byp_alu_rcc_data_e[30]), .A2(byp_alu_rcc_data_e[2]), 
        .A3(byp_alu_rcc_data_e[29]), .A4(byp_alu_rcc_data_e[28]), .Z(n18) );
  HDNOR4D1 U676 ( .A1(byp_alu_rcc_data_e[27]), .A2(byp_alu_rcc_data_e[26]), 
        .A3(byp_alu_rcc_data_e[25]), .A4(byp_alu_rcc_data_e[24]), .Z(n19) );
  HDNAN4D1 U675 ( .A1(n16), .A2(n17), .A3(n18), .A4(n19), .Z(n10) );
  HDNOR4D1 U674 ( .A1(byp_alu_rcc_data_e[23]), .A2(byp_alu_rcc_data_e[22]), 
        .A3(byp_alu_rcc_data_e[21]), .A4(byp_alu_rcc_data_e[20]), .Z(n12) );
  HDNOR4D1 U673 ( .A1(byp_alu_rcc_data_e[1]), .A2(byp_alu_rcc_data_e[19]), 
        .A3(byp_alu_rcc_data_e[18]), .A4(byp_alu_rcc_data_e[17]), .Z(n13) );
  HDNOR4D1 U672 ( .A1(byp_alu_rcc_data_e[16]), .A2(byp_alu_rcc_data_e[15]), 
        .A3(byp_alu_rcc_data_e[14]), .A4(byp_alu_rcc_data_e[13]), .Z(n14) );
  HDNOR4D1 U671 ( .A1(byp_alu_rcc_data_e[12]), .A2(byp_alu_rcc_data_e[11]), 
        .A3(byp_alu_rcc_data_e[10]), .A4(byp_alu_rcc_data_e[0]), .Z(n15) );
  HDNAN4D1 U670 ( .A1(n12), .A2(n13), .A3(n14), .A4(n15), .Z(n11) );
  HDNOR4D1 U669 ( .A1(n8), .A2(n9), .A3(n10), .A4(n11), .Z(exu_ifu_regz_e) );
  HDNAN2D1 U429 ( .A1(n796), .A2(ecl_alu_log_sel_and_e), .Z(n797) );
  HDOAI211D1 U1067 ( .A1(n959), .A2(n796), .B(n965), .C(n797), .Z(n793) );
  HDNOR2D1 U428 ( .A1(byp_alu_rs2_data_e_l[19]), .A2(n422), .Z(n794) );
  HDINVD1 U427 ( .A(byp_alu_rs1_data_e[19]), .Z(n127) );
  HDAOI211D1 U1066 ( .A1(byp_alu_rs1_data_e[19]), .A2(n793), .B(n794), .C(n795), .Z(n197) );
  HDNAN2D1 U417 ( .A1(n782), .A2(ecl_alu_log_sel_and_e), .Z(n783) );
  HDOAI211D1 U1059 ( .A1(n958), .A2(n782), .B(n967), .C(n783), .Z(n779) );
  HDNOR2D1 U416 ( .A1(byp_alu_rs2_data_e_l[20]), .A2(n422), .Z(n780) );
  HDINVD1 U415 ( .A(byp_alu_rs1_data_e[20]), .Z(n129) );
  HDAOI211D1 U1058 ( .A1(byp_alu_rs1_data_e[20]), .A2(n779), .B(n780), .C(n781), .Z(n198) );
  HDNAN2D1 U411 ( .A1(n775), .A2(ecl_alu_log_sel_and_e), .Z(n776) );
  HDOAI211D1 U1055 ( .A1(n957), .A2(n775), .B(n963), .C(n776), .Z(n772) );
  HDNOR2D1 U410 ( .A1(byp_alu_rs2_data_e_l[21]), .A2(n422), .Z(n773) );
  HDINVD1 U409 ( .A(byp_alu_rs1_data_e[21]), .Z(n126) );
  HDAOI211D1 U1054 ( .A1(byp_alu_rs1_data_e[21]), .A2(n772), .B(n773), .C(n774), .Z(n199) );
  HDNAN2D1 U405 ( .A1(n768), .A2(ecl_alu_log_sel_and_e), .Z(n769) );
  HDOAI211D1 U1051 ( .A1(n960), .A2(n768), .B(n964), .C(n769), .Z(n765) );
  HDNOR2D1 U404 ( .A1(byp_alu_rs2_data_e_l[22]), .A2(n422), .Z(n766) );
  HDINVD1 U403 ( .A(byp_alu_rs1_data_e[22]), .Z(n136) );
  HDAOI211D1 U1050 ( .A1(byp_alu_rs1_data_e[22]), .A2(n765), .B(n766), .C(n767), .Z(n200) );
  HDNAN2D1 U453 ( .A1(n824), .A2(ecl_alu_log_sel_and_e), .Z(n825) );
  HDOAI211D1 U1083 ( .A1(n961), .A2(n824), .B(n964), .C(n825), .Z(n821) );
  HDNOR2D1 U452 ( .A1(byp_alu_rs2_data_e_l[15]), .A2(n422), .Z(n822) );
  HDINVD1 U451 ( .A(byp_alu_rs1_data_e[15]), .Z(n121) );
  HDAOI211D1 U1082 ( .A1(byp_alu_rs1_data_e[15]), .A2(n821), .B(n822), .C(n823), .Z(n193) );
  HDNAN2D1 U447 ( .A1(n817), .A2(ecl_alu_log_sel_and_e), .Z(n818) );
  HDOAI211D1 U1079 ( .A1(n958), .A2(n817), .B(n967), .C(n818), .Z(n814) );
  HDNOR2D1 U446 ( .A1(byp_alu_rs2_data_e_l[16]), .A2(n422), .Z(n815) );
  HDINVD1 U445 ( .A(byp_alu_rs1_data_e[16]), .Z(n119) );
  HDAOI211D1 U1078 ( .A1(byp_alu_rs1_data_e[16]), .A2(n814), .B(n815), .C(n816), .Z(n194) );
  HDNAN2D1 U441 ( .A1(n810), .A2(ecl_alu_log_sel_and_e), .Z(n811) );
  HDOAI211D1 U1075 ( .A1(n960), .A2(n810), .B(n965), .C(n811), .Z(n807) );
  HDNOR2D1 U440 ( .A1(byp_alu_rs2_data_e_l[17]), .A2(n422), .Z(n808) );
  HDINVD1 U439 ( .A(byp_alu_rs1_data_e[17]), .Z(n120) );
  HDAOI211D1 U1074 ( .A1(byp_alu_rs1_data_e[17]), .A2(n807), .B(n808), .C(n809), .Z(n195) );
  HDNAN2D1 U435 ( .A1(n803), .A2(ecl_alu_log_sel_and_e), .Z(n804) );
  HDOAI211D1 U1071 ( .A1(n961), .A2(n803), .B(n967), .C(n804), .Z(n800) );
  HDNOR2D1 U434 ( .A1(byp_alu_rs2_data_e_l[18]), .A2(n422), .Z(n801) );
  HDINVD1 U433 ( .A(byp_alu_rs1_data_e[18]), .Z(n128) );
  HDAOI211D1 U1070 ( .A1(byp_alu_rs1_data_e[18]), .A2(n800), .B(n801), .C(n802), .Z(n196) );
  HDNAN2D1 U375 ( .A1(n733), .A2(ecl_alu_log_sel_and_e), .Z(n734) );
  HDOAI211D1 U1031 ( .A1(n957), .A2(n733), .B(n963), .C(n734), .Z(n730) );
  HDNOR2D1 U374 ( .A1(byp_alu_rs2_data_e_l[27]), .A2(n422), .Z(n731) );
  HDINVD1 U373 ( .A(byp_alu_rs1_data_e[27]), .Z(n147) );
  HDAOI211D1 U1030 ( .A1(byp_alu_rs1_data_e[27]), .A2(n730), .B(n731), .C(n732), .Z(n189) );
  HDNAN2D1 U369 ( .A1(n726), .A2(ecl_alu_log_sel_and_e), .Z(n727) );
  HDOAI211D1 U1027 ( .A1(n958), .A2(n726), .B(n963), .C(n727), .Z(n723) );
  HDNOR2D1 U368 ( .A1(byp_alu_rs2_data_e_l[28]), .A2(n422), .Z(n724) );
  HDINVD1 U367 ( .A(byp_alu_rs1_data_e[28]), .Z(n145) );
  HDAOI211D1 U1026 ( .A1(byp_alu_rs1_data_e[28]), .A2(n723), .B(n724), .C(n725), .Z(n190) );
  HDNAN2D1 U363 ( .A1(n719), .A2(ecl_alu_log_sel_and_e), .Z(n720) );
  HDOAI211D1 U1023 ( .A1(n957), .A2(n719), .B(n963), .C(n720), .Z(n716) );
  HDNOR2D1 U362 ( .A1(byp_alu_rs2_data_e_l[29]), .A2(n422), .Z(n717) );
  HDINVD1 U361 ( .A(byp_alu_rs1_data_e[29]), .Z(n146) );
  HDAOI211D1 U1022 ( .A1(byp_alu_rs1_data_e[29]), .A2(n716), .B(n717), .C(n718), .Z(n191) );
  HDNAN2D1 U351 ( .A1(n705), .A2(ecl_alu_log_sel_and_e), .Z(n706) );
  HDOAI211D1 U1015 ( .A1(n957), .A2(n705), .B(n964), .C(n706), .Z(n702) );
  HDNOR2D1 U350 ( .A1(byp_alu_rs2_data_e_l[30]), .A2(n422), .Z(n703) );
  HDINVD1 U349 ( .A(byp_alu_rs1_data_e[30]), .Z(n148) );
  HDAOI211D1 U1014 ( .A1(byp_alu_rs1_data_e[30]), .A2(n702), .B(n703), .C(n704), .Z(n192) );
  HDNAN2D1 U399 ( .A1(n761), .A2(ecl_alu_log_sel_and_e), .Z(n762) );
  HDOAI211D1 U1047 ( .A1(n960), .A2(n761), .B(n963), .C(n762), .Z(n758) );
  HDNOR2D1 U398 ( .A1(byp_alu_rs2_data_e_l[23]), .A2(n422), .Z(n759) );
  HDINVD1 U397 ( .A(byp_alu_rs1_data_e[23]), .Z(n135) );
  HDAOI211D1 U1046 ( .A1(byp_alu_rs1_data_e[23]), .A2(n758), .B(n759), .C(n760), .Z(n185) );
  HDNAN2D1 U393 ( .A1(n754), .A2(ecl_alu_log_sel_and_e), .Z(n755) );
  HDOAI211D1 U1043 ( .A1(n961), .A2(n754), .B(n963), .C(n755), .Z(n751) );
  HDNOR2D1 U392 ( .A1(byp_alu_rs2_data_e_l[24]), .A2(n422), .Z(n752) );
  HDINVD1 U391 ( .A(byp_alu_rs1_data_e[24]), .Z(n137) );
  HDAOI211D1 U1042 ( .A1(byp_alu_rs1_data_e[24]), .A2(n751), .B(n752), .C(n753), .Z(n186) );
  HDNAN2D1 U387 ( .A1(n747), .A2(ecl_alu_log_sel_and_e), .Z(n748) );
  HDOAI211D1 U1039 ( .A1(n962), .A2(n747), .B(n963), .C(n748), .Z(n744) );
  HDNOR2D1 U386 ( .A1(byp_alu_rs2_data_e_l[25]), .A2(n422), .Z(n745) );
  HDINVD1 U385 ( .A(byp_alu_rs1_data_e[25]), .Z(n138) );
  HDAOI211D1 U1038 ( .A1(byp_alu_rs1_data_e[25]), .A2(n744), .B(n745), .C(n746), .Z(n187) );
  HDNAN2D1 U381 ( .A1(n740), .A2(ecl_alu_log_sel_and_e), .Z(n741) );
  HDOAI211D1 U1035 ( .A1(n959), .A2(n740), .B(n963), .C(n741), .Z(n737) );
  HDNOR2D1 U380 ( .A1(byp_alu_rs2_data_e_l[26]), .A2(n422), .Z(n738) );
  HDINVD1 U379 ( .A(byp_alu_rs1_data_e[26]), .Z(n134) );
  HDAOI211D1 U1034 ( .A1(byp_alu_rs1_data_e[26]), .A2(n737), .B(n738), .C(n739), .Z(n188) );
  HDNOR4D1 U756 ( .A1(n181), .A2(n182), .A3(n183), .A4(n184), .Z(n28) );
  HDNAN2D1 U291 ( .A1(n635), .A2(ecl_alu_log_sel_and_e), .Z(n636) );
  HDOAI211D1 U973 ( .A1(n958), .A2(n635), .B(n965), .C(n636), .Z(n632) );
  HDNOR2D1 U290 ( .A1(byp_alu_rs2_data_e_l[3]), .A2(n422), .Z(n633) );
  HDINVD1 U289 ( .A(byp_alu_rs1_data_e[3]), .Z(n85) );
  HDAOI211D1 U972 ( .A1(byp_alu_rs1_data_e[3]), .A2(n632), .B(n633), .C(n634), 
        .Z(n177) );
  HDNAN2D1 U225 ( .A1(n558), .A2(ecl_alu_log_sel_and_e), .Z(n559) );
  HDOAI211D1 U929 ( .A1(n960), .A2(n558), .B(n967), .C(n559), .Z(n555) );
  HDNOR2D1 U224 ( .A1(byp_alu_rs2_data_e_l[4]), .A2(n422), .Z(n556) );
  HDINVD1 U223 ( .A(byp_alu_rs1_data_e[4]), .Z(n160) );
  HDAOI211D1 U928 ( .A1(byp_alu_rs1_data_e[4]), .A2(n555), .B(n556), .C(n557), 
        .Z(n178) );
  HDNAN2D1 U159 ( .A1(n481), .A2(ecl_alu_log_sel_and_e), .Z(n482) );
  HDOAI211D1 U885 ( .A1(n961), .A2(n481), .B(n968), .C(n482), .Z(n478) );
  HDNOR2D1 U158 ( .A1(byp_alu_rs2_data_e_l[5]), .A2(n422), .Z(n479) );
  HDINVD1 U157 ( .A(byp_alu_rs1_data_e[5]), .Z(n157) );
  HDAOI211D1 U884 ( .A1(byp_alu_rs1_data_e[5]), .A2(n478), .B(n479), .C(n480), 
        .Z(n179) );
  HDNAN2D1 U129 ( .A1(n446), .A2(ecl_alu_log_sel_and_e), .Z(n447) );
  HDOAI211D1 U865 ( .A1(n962), .A2(n446), .B(n966), .C(n447), .Z(n443) );
  HDNOR2D1 U128 ( .A1(byp_alu_rs2_data_e_l[6]), .A2(n422), .Z(n444) );
  HDINVD1 U127 ( .A(byp_alu_rs1_data_e[6]), .Z(n159) );
  HDAOI211D1 U864 ( .A1(byp_alu_rs1_data_e[6]), .A2(n443), .B(n444), .C(n445), 
        .Z(n180) );
  HDINVD1 U345 ( .A(byp_alu_rs1_data_e[31]), .Z(n143) );
  HDAOI32D1 U1011 ( .A1(ecl_alu_log_sel_xor_e), .A2(n698), .A3(n143), .B1(
        ecl_alu_log_sel_or_e), .B2(n698), .Z(n695) );
  HDNAN2D1 U344 ( .A1(n698), .A2(ecl_alu_log_sel_and_e), .Z(n699) );
  HDOAI211D1 U1010 ( .A1(n957), .A2(n698), .B(n964), .C(n699), .Z(n697) );
  HDNAN2D1 U343 ( .A1(byp_alu_rs1_data_e[31]), .A2(n697), .Z(n696) );
  HDOAI211D1 U1009 ( .A1(byp_alu_rs2_data_e_l[31]), .A2(n422), .B(n695), .C(
        n696), .Z(alu_ecl_log_n32_e) );
  HDINVD1 U342 ( .A(alu_ecl_log_n32_e), .Z(n173) );
  HDNAN2D1 U493 ( .A1(n866), .A2(ecl_alu_log_sel_and_e), .Z(n867) );
  HDOAI211D1 U1107 ( .A1(n958), .A2(n866), .B(n966), .C(n867), .Z(n863) );
  HDNOR2D1 U491 ( .A1(byp_alu_rs2_data_e_l[0]), .A2(n422), .Z(n864) );
  HDINVD1 U490 ( .A(byp_alu_rs1_data_e[0]), .Z(n86) );
  HDAOI211D1 U1106 ( .A1(byp_alu_rs1_data_e[0]), .A2(n863), .B(n864), .C(n865), 
        .Z(n174) );
  HDNAN2D1 U423 ( .A1(n789), .A2(ecl_alu_log_sel_and_e), .Z(n790) );
  HDOAI211D1 U1063 ( .A1(n962), .A2(n789), .B(n968), .C(n790), .Z(n786) );
  HDNOR2D1 U422 ( .A1(byp_alu_rs2_data_e_l[1]), .A2(n422), .Z(n787) );
  HDINVD1 U421 ( .A(byp_alu_rs1_data_e[1]), .Z(n80) );
  HDAOI211D1 U1062 ( .A1(byp_alu_rs1_data_e[1]), .A2(n786), .B(n787), .C(n788), 
        .Z(n175) );
  HDNAN2D1 U357 ( .A1(n712), .A2(ecl_alu_log_sel_and_e), .Z(n713) );
  HDOAI211D1 U1019 ( .A1(n957), .A2(n712), .B(n964), .C(n713), .Z(n709) );
  HDNOR2D1 U356 ( .A1(byp_alu_rs2_data_e_l[2]), .A2(n422), .Z(n710) );
  HDINVD1 U355 ( .A(byp_alu_rs1_data_e[2]), .Z(n81) );
  HDAOI211D1 U1018 ( .A1(byp_alu_rs1_data_e[2]), .A2(n709), .B(n710), .C(n711), 
        .Z(n176) );
  HDNAN2D1 U477 ( .A1(n852), .A2(ecl_alu_log_sel_and_e), .Z(n853) );
  HDOAI211D1 U1099 ( .A1(n960), .A2(n852), .B(n965), .C(n853), .Z(n849) );
  HDNOR2D1 U476 ( .A1(byp_alu_rs2_data_e_l[11]), .A2(n422), .Z(n850) );
  HDINVD1 U475 ( .A(byp_alu_rs1_data_e[11]), .Z(n110) );
  HDAOI211D1 U1098 ( .A1(byp_alu_rs1_data_e[11]), .A2(n849), .B(n850), .C(n851), .Z(n169) );
  HDNAN2D1 U471 ( .A1(n845), .A2(ecl_alu_log_sel_and_e), .Z(n846) );
  HDOAI211D1 U1095 ( .A1(n961), .A2(n845), .B(n964), .C(n846), .Z(n842) );
  HDNOR2D1 U470 ( .A1(byp_alu_rs2_data_e_l[12]), .A2(n422), .Z(n843) );
  HDINVD1 U469 ( .A(byp_alu_rs1_data_e[12]), .Z(n153) );
  HDAOI211D1 U1094 ( .A1(byp_alu_rs1_data_e[12]), .A2(n842), .B(n843), .C(n844), .Z(n170) );
  HDNAN2D1 U465 ( .A1(n838), .A2(ecl_alu_log_sel_and_e), .Z(n839) );
  HDOAI211D1 U1091 ( .A1(n962), .A2(n838), .B(n968), .C(n839), .Z(n835) );
  HDNOR2D1 U464 ( .A1(byp_alu_rs2_data_e_l[13]), .A2(n422), .Z(n836) );
  HDINVD1 U463 ( .A(byp_alu_rs1_data_e[13]), .Z(n107) );
  HDAOI211D1 U1090 ( .A1(byp_alu_rs1_data_e[13]), .A2(n835), .B(n836), .C(n837), .Z(n171) );
  HDNAN2D1 U459 ( .A1(n831), .A2(ecl_alu_log_sel_and_e), .Z(n832) );
  HDOAI211D1 U1087 ( .A1(n959), .A2(n831), .B(n966), .C(n832), .Z(n828) );
  HDNOR2D1 U458 ( .A1(byp_alu_rs2_data_e_l[14]), .A2(n422), .Z(n829) );
  HDINVD1 U457 ( .A(byp_alu_rs1_data_e[14]), .Z(n108) );
  HDAOI211D1 U1086 ( .A1(byp_alu_rs1_data_e[14]), .A2(n828), .B(n829), .C(n830), .Z(n172) );
  HDNAN2D1 U123 ( .A1(n439), .A2(ecl_alu_log_sel_and_e), .Z(n440) );
  HDOAI211D1 U861 ( .A1(n962), .A2(n439), .B(n963), .C(n440), .Z(n436) );
  HDNOR2D1 U122 ( .A1(byp_alu_rs2_data_e_l[7]), .A2(n422), .Z(n437) );
  HDINVD1 U121 ( .A(byp_alu_rs1_data_e[7]), .Z(n155) );
  HDAOI211D1 U860 ( .A1(byp_alu_rs1_data_e[7]), .A2(n436), .B(n437), .C(n438), 
        .Z(n165) );
  HDNAN2D1 U117 ( .A1(n432), .A2(ecl_alu_log_sel_and_e), .Z(n433) );
  HDOAI211D1 U857 ( .A1(n962), .A2(n432), .B(n964), .C(n433), .Z(n429) );
  HDNOR2D1 U116 ( .A1(byp_alu_rs2_data_e_l[8]), .A2(n422), .Z(n430) );
  HDINVD1 U115 ( .A(byp_alu_rs1_data_e[8]), .Z(n156) );
  HDAOI211D1 U856 ( .A1(byp_alu_rs1_data_e[8]), .A2(n429), .B(n430), .C(n431), 
        .Z(n166) );
  HDNAN2D1 U111 ( .A1(n421), .A2(ecl_alu_log_sel_and_e), .Z(n425) );
  HDOAI211D1 U853 ( .A1(n962), .A2(n421), .B(n965), .C(n425), .Z(n418) );
  HDNOR2D1 U110 ( .A1(byp_alu_rs2_data_e_l[9]), .A2(n422), .Z(n419) );
  HDINVD1 U109 ( .A(byp_alu_rs1_data_e[9]), .Z(n158) );
  HDAOI211D1 U852 ( .A1(byp_alu_rs1_data_e[9]), .A2(n418), .B(n419), .C(n420), 
        .Z(n167) );
  HDNAN2D1 U483 ( .A1(n859), .A2(ecl_alu_log_sel_and_e), .Z(n860) );
  HDOAI211D1 U1103 ( .A1(n957), .A2(n859), .B(n963), .C(n860), .Z(n856) );
  HDNOR2D1 U482 ( .A1(byp_alu_rs2_data_e_l[10]), .A2(n422), .Z(n857) );
  HDINVD1 U481 ( .A(byp_alu_rs1_data_e[10]), .Z(n154) );
  HDAOI211D1 U1102 ( .A1(byp_alu_rs1_data_e[10]), .A2(n856), .B(n857), .C(n858), .Z(n168) );
  HDNOR4D1 U751 ( .A1(n161), .A2(n162), .A3(n163), .A4(n164), .Z(n29) );
  HDNOR4D1 U746 ( .A1(n149), .A2(n150), .A3(n151), .A4(n152), .Z(n53) );
  HDINVD1 U46 ( .A(alu_ecl_adderin2_31_e), .Z(n144) );
  HDNAN4D1 U741 ( .A1(n139), .A2(n140), .A3(n141), .A4(n142), .Z(n111) );
  HDAOI22D1 U737 ( .A1(byp_alu_rs1_data_e[23]), .A2(n96), .B1(
        byp_alu_rs1_data_e[24]), .B2(n92), .Z(n133) );
  HDNAN4D1 U736 ( .A1(n130), .A2(n131), .A3(n132), .A4(n133), .Z(n112) );
  HDAOI22D1 U734 ( .A1(byp_alu_rs1_data_e[17]), .A2(n106), .B1(
        byp_alu_rs1_data_e[18]), .B2(n98), .Z(n123) );
  HDNAN4D1 U731 ( .A1(n122), .A2(n123), .A3(n124), .A4(n125), .Z(n113) );
  HDNAN4D1 U726 ( .A1(n115), .A2(n116), .A3(n117), .A4(n118), .Z(n114) );
  HDOR4D1 U725 ( .A1(n111), .A2(n112), .A3(n113), .A4(n114), .Z(n73) );
  HDNOR4D1 U720 ( .A1(n99), .A2(n100), .A3(n101), .A4(n102), .Z(n75) );
  HDNOR4D1 U715 ( .A1(n87), .A2(n88), .A3(n89), .A4(n90), .Z(n76) );
  HDNAN2D1 U10 ( .A1(addsub_rs2_data_0), .A2(n82), .Z(n83) );
  HDOAI211D1 U713 ( .A1(n82), .A2(addsub_rs2_data_0), .B(n83), .C(n84), .Z(n78) );
  HDAOI211D1 U711 ( .A1(n60), .A2(byp_alu_rs1_data_e[30]), .B(n78), .C(n79), 
        .Z(n77) );
  HDNAN3D1 U6 ( .A1(n75), .A2(n76), .A3(n77), .Z(n74) );
  HDAOI211D1 U710 ( .A1(byp_alu_rs1_data_e[29]), .A2(n63), .B(n73), .C(n74), 
        .Z(n54) );
  HDOR2D1 U709 ( .A1(addsub_rs2_data_0), .A2(byp_alu_rs1_data_e[0]), .Z(n72)
         );
  HDAOI22D1 U705 ( .A1(byp_alu_rs1_data_e[11]), .A2(n70), .B1(
        byp_alu_rs1_data_e[13]), .B2(n69), .Z(n66) );
  HDNAN4D1 U703 ( .A1(n64), .A2(n65), .A3(n66), .A4(n67), .Z(n57) );
  HDNOR3D1 U5 ( .A1(n57), .A2(n58), .A3(n59), .Z(n56) );
  HDNAN4D1 U700 ( .A1(n53), .A2(n54), .A3(n55), .A4(n56), .Z(n32) );
  HDAOI22D1 U699 ( .A1(byp_alu_rs1_data_e[1]), .A2(n52), .B1(
        byp_alu_rs1_data_e[3]), .B2(n51), .Z(n45) );
  HDAOI22D1 U696 ( .A1(byp_alu_rs1_data_e[4]), .A2(n49), .B1(
        byp_alu_rs1_data_e[6]), .B2(n44), .Z(n48) );
  HDNAN4D1 U695 ( .A1(n45), .A2(n46), .A3(n47), .A4(n48), .Z(n33) );
  HDAOI22D1 U691 ( .A1(byp_alu_rs1_data_e[8]), .A2(n39), .B1(
        byp_alu_rs1_data_e[10]), .B2(n40), .Z(n38) );
  HDNAN4D1 U690 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .Z(n34) );
  HDNOR3D1 U4 ( .A1(n32), .A2(n33), .A3(n34), .Z(n31) );
  HDNAN2D1 U213 ( .A1(n544), .A2(ecl_alu_log_sel_and_e), .Z(n545) );
  HDOAI211D1 U921 ( .A1(n960), .A2(n544), .B(n967), .C(n545), .Z(n541) );
  HDNOR2D1 U212 ( .A1(byp_alu_rs2_data_e_l[51]), .A2(n450), .Z(n542) );
  HDINVD1 U211 ( .A(byp_alu_rs1_data_e[51]), .Z(n282) );
  HDAOI211D1 U920 ( .A1(byp_alu_rs1_data_e[51]), .A2(n541), .B(n542), .C(n543), 
        .Z(n370) );
  HDNAN2D1 U207 ( .A1(n537), .A2(ecl_alu_log_sel_and_e), .Z(n538) );
  HDOAI211D1 U917 ( .A1(n960), .A2(n537), .B(n967), .C(n538), .Z(n534) );
  HDNOR2D1 U206 ( .A1(byp_alu_rs2_data_e_l[52]), .A2(n450), .Z(n535) );
  HDINVD1 U205 ( .A(byp_alu_rs1_data_e[52]), .Z(n284) );
  HDAOI211D1 U916 ( .A1(byp_alu_rs1_data_e[52]), .A2(n534), .B(n535), .C(n536), 
        .Z(n371) );
  HDNAN2D1 U201 ( .A1(n530), .A2(ecl_alu_log_sel_and_e), .Z(n531) );
  HDOAI211D1 U913 ( .A1(n960), .A2(n530), .B(n967), .C(n531), .Z(n527) );
  HDINVD1 U199 ( .A(byp_alu_rs1_data_e[53]), .Z(n280) );
  HDAOI211D1 U912 ( .A1(byp_alu_rs1_data_e[53]), .A2(n527), .B(n528), .C(n529), 
        .Z(n372) );
  HDNAN2D1 U195 ( .A1(n523), .A2(ecl_alu_log_sel_and_e), .Z(n524) );
  HDOAI211D1 U909 ( .A1(n961), .A2(n523), .B(n967), .C(n524), .Z(n520) );
  HDINVD1 U193 ( .A(byp_alu_rs1_data_e[54]), .Z(n281) );
  HDAOI211D1 U908 ( .A1(byp_alu_rs1_data_e[54]), .A2(n520), .B(n521), .C(n522), 
        .Z(n373) );
  HDNAN2D1 U243 ( .A1(n579), .A2(ecl_alu_log_sel_and_e), .Z(n580) );
  HDOAI211D1 U941 ( .A1(n959), .A2(n579), .B(n966), .C(n580), .Z(n576) );
  HDINVD1 U241 ( .A(byp_alu_rs1_data_e[47]), .Z(n311) );
  HDAOI211D1 U940 ( .A1(byp_alu_rs1_data_e[47]), .A2(n576), .B(n577), .C(n578), 
        .Z(n366) );
  HDNAN2D1 U237 ( .A1(n572), .A2(ecl_alu_log_sel_and_e), .Z(n573) );
  HDOAI211D1 U937 ( .A1(n960), .A2(n572), .B(n966), .C(n573), .Z(n569) );
  HDNOR2D1 U236 ( .A1(byp_alu_rs2_data_e_l[48]), .A2(n941), .Z(n570) );
  HDINVD1 U235 ( .A(byp_alu_rs1_data_e[48]), .Z(n309) );
  HDAOI211D1 U936 ( .A1(byp_alu_rs1_data_e[48]), .A2(n569), .B(n570), .C(n571), 
        .Z(n367) );
  HDNAN2D1 U231 ( .A1(n565), .A2(ecl_alu_log_sel_and_e), .Z(n566) );
  HDOAI211D1 U933 ( .A1(n960), .A2(n565), .B(n967), .C(n566), .Z(n562) );
  HDINVD1 U229 ( .A(byp_alu_rs1_data_e[49]), .Z(n291) );
  HDAOI211D1 U932 ( .A1(byp_alu_rs1_data_e[49]), .A2(n562), .B(n563), .C(n564), 
        .Z(n368) );
  HDNAN2D1 U219 ( .A1(n551), .A2(ecl_alu_log_sel_and_e), .Z(n552) );
  HDOAI211D1 U925 ( .A1(n960), .A2(n551), .B(n967), .C(n552), .Z(n548) );
  HDINVD1 U217 ( .A(byp_alu_rs1_data_e[50]), .Z(n285) );
  HDAOI211D1 U924 ( .A1(byp_alu_rs1_data_e[50]), .A2(n548), .B(n549), .C(n550), 
        .Z(n369) );
  HDNAN2D1 U165 ( .A1(n488), .A2(ecl_alu_log_sel_and_e), .Z(n489) );
  HDOAI211D1 U889 ( .A1(n961), .A2(n488), .B(n968), .C(n489), .Z(n485) );
  HDNOR2D1 U164 ( .A1(byp_alu_rs2_data_e_l[59]), .A2(n450), .Z(n486) );
  HDINVD1 U163 ( .A(byp_alu_rs1_data_e[59]), .Z(n265) );
  HDAOI211D1 U888 ( .A1(byp_alu_rs1_data_e[59]), .A2(n485), .B(n486), .C(n487), 
        .Z(n362) );
  HDNAN2D1 U153 ( .A1(n474), .A2(ecl_alu_log_sel_and_e), .Z(n475) );
  HDOAI211D1 U881 ( .A1(n962), .A2(n474), .B(n968), .C(n475), .Z(n471) );
  HDNOR2D1 U152 ( .A1(byp_alu_rs2_data_e_l[60]), .A2(n450), .Z(n472) );
  HDINVD1 U151 ( .A(byp_alu_rs1_data_e[60]), .Z(n266) );
  HDAOI211D1 U880 ( .A1(byp_alu_rs1_data_e[60]), .A2(n471), .B(n472), .C(n473), 
        .Z(n363) );
  HDNAN2D1 U147 ( .A1(n467), .A2(ecl_alu_log_sel_and_e), .Z(n468) );
  HDOAI211D1 U877 ( .A1(n962), .A2(n467), .B(n967), .C(n468), .Z(n464) );
  HDNOR2D1 U146 ( .A1(byp_alu_rs2_data_e_l[61]), .A2(n450), .Z(n465) );
  HDINVD1 U145 ( .A(byp_alu_rs1_data_e[61]), .Z(n268) );
  HDAOI211D1 U876 ( .A1(byp_alu_rs1_data_e[61]), .A2(n464), .B(n465), .C(n466), 
        .Z(n364) );
  HDNAN2D1 U141 ( .A1(n460), .A2(ecl_alu_log_sel_and_e), .Z(n461) );
  HDOAI211D1 U873 ( .A1(n962), .A2(n460), .B(n968), .C(n461), .Z(n457) );
  HDNOR2D1 U140 ( .A1(byp_alu_rs2_data_e_l[62]), .A2(n450), .Z(n458) );
  HDINVD1 U139 ( .A(byp_alu_rs1_data_e[62]), .Z(n270) );
  HDAOI211D1 U872 ( .A1(byp_alu_rs1_data_e[62]), .A2(n457), .B(n458), .C(n459), 
        .Z(n365) );
  HDNAN2D1 U189 ( .A1(n516), .A2(ecl_alu_log_sel_and_e), .Z(n517) );
  HDOAI211D1 U905 ( .A1(n961), .A2(n516), .B(n968), .C(n517), .Z(n513) );
  HDINVD1 U187 ( .A(byp_alu_rs1_data_e[55]), .Z(n283) );
  HDAOI211D1 U904 ( .A1(byp_alu_rs1_data_e[55]), .A2(n513), .B(n514), .C(n515), 
        .Z(n358) );
  HDNAN2D1 U183 ( .A1(n509), .A2(ecl_alu_log_sel_and_e), .Z(n510) );
  HDOAI211D1 U901 ( .A1(n961), .A2(n509), .B(n968), .C(n510), .Z(n506) );
  HDINVD1 U181 ( .A(byp_alu_rs1_data_e[56]), .Z(n275) );
  HDAOI211D1 U900 ( .A1(byp_alu_rs1_data_e[56]), .A2(n506), .B(n507), .C(n508), 
        .Z(n359) );
  HDNAN2D1 U177 ( .A1(n502), .A2(ecl_alu_log_sel_and_e), .Z(n503) );
  HDOAI211D1 U897 ( .A1(n961), .A2(n502), .B(n968), .C(n503), .Z(n499) );
  HDINVD1 U175 ( .A(byp_alu_rs1_data_e[57]), .Z(n267) );
  HDAOI211D1 U896 ( .A1(byp_alu_rs1_data_e[57]), .A2(n499), .B(n500), .C(n501), 
        .Z(n360) );
  HDNAN2D1 U171 ( .A1(n495), .A2(ecl_alu_log_sel_and_e), .Z(n496) );
  HDOAI211D1 U893 ( .A1(n961), .A2(n495), .B(n968), .C(n496), .Z(n492) );
  HDINVD1 U169 ( .A(byp_alu_rs1_data_e[58]), .Z(n271) );
  HDAOI211D1 U892 ( .A1(byp_alu_rs1_data_e[58]), .A2(n492), .B(n493), .C(n494), 
        .Z(n361) );
  HDNOR4D1 U831 ( .A1(n354), .A2(n355), .A3(n356), .A4(n357), .Z(n201) );
  HDNAN2D1 U321 ( .A1(n670), .A2(ecl_alu_log_sel_and_e), .Z(n671) );
  HDOAI211D1 U993 ( .A1(n958), .A2(n670), .B(n964), .C(n671), .Z(n667) );
  HDINVD1 U319 ( .A(byp_alu_rs1_data_e[35]), .Z(n333) );
  HDAOI211D1 U992 ( .A1(byp_alu_rs1_data_e[35]), .A2(n667), .B(n668), .C(n669), 
        .Z(n350) );
  HDNAN2D1 U315 ( .A1(n663), .A2(ecl_alu_log_sel_and_e), .Z(n664) );
  HDOAI211D1 U989 ( .A1(n958), .A2(n663), .B(n965), .C(n664), .Z(n660) );
  HDINVD1 U313 ( .A(byp_alu_rs1_data_e[36]), .Z(n332) );
  HDAOI211D1 U988 ( .A1(byp_alu_rs1_data_e[36]), .A2(n660), .B(n661), .C(n662), 
        .Z(n351) );
  HDNAN2D1 U309 ( .A1(n656), .A2(ecl_alu_log_sel_and_e), .Z(n657) );
  HDOAI211D1 U985 ( .A1(n958), .A2(n656), .B(n965), .C(n657), .Z(n653) );
  HDINVD1 U307 ( .A(byp_alu_rs1_data_e[37]), .Z(n331) );
  HDAOI211D1 U984 ( .A1(byp_alu_rs1_data_e[37]), .A2(n653), .B(n654), .C(n655), 
        .Z(n352) );
  HDNAN2D1 U303 ( .A1(n649), .A2(ecl_alu_log_sel_and_e), .Z(n650) );
  HDOAI211D1 U981 ( .A1(n958), .A2(n649), .B(n965), .C(n650), .Z(n646) );
  HDINVD1 U301 ( .A(byp_alu_rs1_data_e[38]), .Z(n330) );
  HDAOI211D1 U980 ( .A1(byp_alu_rs1_data_e[38]), .A2(n646), .B(n647), .C(n648), 
        .Z(n353) );
  HDINVD1 U133 ( .A(byp_alu_rs1_data_e[63]), .Z(n304) );
  HDAOI32D1 U869 ( .A1(n453), .A2(n304), .A3(ecl_alu_log_sel_xor_e), .B1(
        ecl_alu_log_sel_or_e), .B2(n453), .Z(n452) );
  HDOAI211D1 U868 ( .A1(byp_alu_rs2_data_e_l[63]), .A2(n450), .B(n451), .C(
        n452), .Z(alu_ecl_log_n64_e) );
  HDINVD1 U132 ( .A(alu_ecl_log_n64_e), .Z(n346) );
  HDNAN2D1 U339 ( .A1(n691), .A2(ecl_alu_log_sel_and_e), .Z(n692) );
  HDOAI211D1 U1006 ( .A1(n957), .A2(n691), .B(n964), .C(n692), .Z(n688) );
  HDINVD1 U337 ( .A(byp_alu_rs1_data_e[32]), .Z(n315) );
  HDAOI211D1 U1004 ( .A1(byp_alu_rs1_data_e[32]), .A2(n688), .B(n689), .C(n690), .Z(n347) );
  HDNAN2D1 U333 ( .A1(n684), .A2(ecl_alu_log_sel_and_e), .Z(n685) );
  HDOAI211D1 U1001 ( .A1(n957), .A2(n684), .B(n964), .C(n685), .Z(n681) );
  HDNOR2D1 U332 ( .A1(byp_alu_rs2_data_e_l[33]), .A2(n450), .Z(n682) );
  HDINVD1 U331 ( .A(byp_alu_rs1_data_e[33]), .Z(n314) );
  HDAOI211D1 U1000 ( .A1(byp_alu_rs1_data_e[33]), .A2(n681), .B(n682), .C(n683), .Z(n348) );
  HDNAN2D1 U327 ( .A1(n677), .A2(ecl_alu_log_sel_and_e), .Z(n678) );
  HDOAI211D1 U997 ( .A1(n957), .A2(n677), .B(n964), .C(n678), .Z(n674) );
  HDINVD1 U325 ( .A(byp_alu_rs1_data_e[34]), .Z(n313) );
  HDAOI211D1 U996 ( .A1(byp_alu_rs1_data_e[34]), .A2(n674), .B(n675), .C(n676), 
        .Z(n349) );
  HDNAN2D1 U267 ( .A1(n607), .A2(ecl_alu_log_sel_and_e), .Z(n608) );
  HDOAI211D1 U957 ( .A1(n959), .A2(n607), .B(n966), .C(n608), .Z(n604) );
  HDINVD1 U265 ( .A(byp_alu_rs1_data_e[43]), .Z(n321) );
  HDAOI211D1 U956 ( .A1(byp_alu_rs1_data_e[43]), .A2(n604), .B(n605), .C(n606), 
        .Z(n342) );
  HDNAN2D1 U261 ( .A1(n600), .A2(ecl_alu_log_sel_and_e), .Z(n601) );
  HDOAI211D1 U953 ( .A1(n959), .A2(n600), .B(n966), .C(n601), .Z(n597) );
  HDINVD1 U259 ( .A(byp_alu_rs1_data_e[44]), .Z(n320) );
  HDAOI211D1 U952 ( .A1(byp_alu_rs1_data_e[44]), .A2(n597), .B(n598), .C(n599), 
        .Z(n343) );
  HDNAN2D1 U255 ( .A1(n593), .A2(ecl_alu_log_sel_and_e), .Z(n594) );
  HDOAI211D1 U949 ( .A1(n959), .A2(n593), .B(n966), .C(n594), .Z(n590) );
  HDINVD1 U253 ( .A(byp_alu_rs1_data_e[45]), .Z(n312) );
  HDAOI211D1 U948 ( .A1(byp_alu_rs1_data_e[45]), .A2(n590), .B(n591), .C(n592), 
        .Z(n344) );
  HDNAN2D1 U249 ( .A1(n586), .A2(ecl_alu_log_sel_and_e), .Z(n587) );
  HDOAI211D1 U945 ( .A1(n959), .A2(n586), .B(n966), .C(n587), .Z(n583) );
  HDINVD1 U247 ( .A(byp_alu_rs1_data_e[46]), .Z(n310) );
  HDAOI211D1 U944 ( .A1(byp_alu_rs1_data_e[46]), .A2(n583), .B(n584), .C(n585), 
        .Z(n345) );
  HDNAN2D1 U297 ( .A1(n642), .A2(ecl_alu_log_sel_and_e), .Z(n643) );
  HDOAI211D1 U977 ( .A1(n958), .A2(n642), .B(n965), .C(n643), .Z(n639) );
  HDINVD1 U295 ( .A(byp_alu_rs1_data_e[39]), .Z(n329) );
  HDAOI211D1 U976 ( .A1(byp_alu_rs1_data_e[39]), .A2(n639), .B(n640), .C(n641), 
        .Z(n338) );
  HDNAN2D1 U285 ( .A1(n628), .A2(ecl_alu_log_sel_and_e), .Z(n629) );
  HDOAI211D1 U969 ( .A1(n958), .A2(n628), .B(n965), .C(n629), .Z(n625) );
  HDINVD1 U283 ( .A(byp_alu_rs1_data_e[40]), .Z(n324) );
  HDAOI211D1 U968 ( .A1(byp_alu_rs1_data_e[40]), .A2(n625), .B(n626), .C(n627), 
        .Z(n339) );
  HDNAN2D1 U279 ( .A1(n621), .A2(ecl_alu_log_sel_and_e), .Z(n622) );
  HDOAI211D1 U965 ( .A1(n959), .A2(n621), .B(n965), .C(n622), .Z(n618) );
  HDINVD1 U277 ( .A(byp_alu_rs1_data_e[41]), .Z(n323) );
  HDAOI211D1 U964 ( .A1(byp_alu_rs1_data_e[41]), .A2(n618), .B(n619), .C(n620), 
        .Z(n340) );
  HDNAN2D1 U273 ( .A1(n614), .A2(ecl_alu_log_sel_and_e), .Z(n615) );
  HDOAI211D1 U961 ( .A1(n959), .A2(n614), .B(n966), .C(n615), .Z(n611) );
  HDINVD1 U271 ( .A(byp_alu_rs1_data_e[42]), .Z(n322) );
  HDAOI211D1 U960 ( .A1(byp_alu_rs1_data_e[42]), .A2(n611), .B(n612), .C(n613), 
        .Z(n341) );
  HDNOR4D1 U826 ( .A1(n334), .A2(n335), .A3(n336), .A4(n337), .Z(n202) );
  HDAOI22D1 U823 ( .A1(byp_alu_rs1_data_e[36]), .A2(n220), .B1(
        byp_alu_rs1_data_e[38]), .B2(n297), .Z(n327) );
  HDNAN4D1 U821 ( .A1(n325), .A2(n326), .A3(n327), .A4(n328), .Z(n204) );
  HDAOI22D1 U819 ( .A1(byp_alu_rs1_data_e[39]), .A2(n217), .B1(
        byp_alu_rs1_data_e[41]), .B2(n294), .Z(n317) );
  HDNAN4D1 U816 ( .A1(n316), .A2(n317), .A3(n318), .A4(n319), .Z(n205) );
  HDAOI22D1 U808 ( .A1(n218), .A2(byp_alu_rs1_data_e[35]), .B1(n223), .B2(
        byp_alu_rs1_data_e[33]), .Z(n303) );
  HDAOI211D1 U806 ( .A1(n221), .A2(byp_alu_rs1_data_e[32]), .B(n301), .C(n302), 
        .Z(n300) );
  HDNAN3D1 U57 ( .A1(n298), .A2(n299), .A3(n300), .Z(n206) );
  HDNOR4D1 U801 ( .A1(n286), .A2(n287), .A3(n288), .A4(n289), .Z(n272) );
  HDNOR4D1 U796 ( .A1(n276), .A2(n277), .A3(n278), .A4(n279), .Z(n273) );
  HDAND3D1 U794 ( .A1(n272), .A2(n273), .A3(n274), .Z(n208) );
  HDNAN4D1 U784 ( .A1(n254), .A2(n255), .A3(n256), .A4(n257), .Z(n224) );
  HDAOI22D1 U780 ( .A1(byp_alu_rs1_data_e[48]), .A2(n249), .B1(
        byp_alu_rs1_data_e[49]), .B2(n250), .Z(n248) );
  HDNAN4D1 U779 ( .A1(n245), .A2(n246), .A3(n247), .A4(n248), .Z(n225) );
  HDAOI22D1 U775 ( .A1(byp_alu_rs1_data_e[60]), .A2(n242), .B1(
        byp_alu_rs1_data_e[61]), .B2(n243), .Z(n241) );
  HDNAN4D1 U774 ( .A1(n238), .A2(n239), .A3(n240), .A4(n241), .Z(n226) );
  HDAOI22D1 U772 ( .A1(byp_alu_rs1_data_e[54]), .A2(n235), .B1(
        byp_alu_rs1_data_e[55]), .B2(n236), .Z(n229) );
  HDNAN4D1 U769 ( .A1(n228), .A2(n229), .A3(n230), .A4(n231), .Z(n227) );
  HDNOR4D1 U768 ( .A1(n224), .A2(n225), .A3(n226), .A4(n227), .Z(n210) );
  HDNOR4D1 U763 ( .A1(n212), .A2(n213), .A3(n214), .A4(n215), .Z(n211) );
  HDNAN4D1 U762 ( .A1(n208), .A2(n209), .A3(n210), .A4(n211), .Z(n207) );
  HDNOR4D1 U761 ( .A1(n204), .A2(n205), .A3(n206), .A4(n207), .Z(n203) );
  HDMUX2D1 U668 ( .A0(exu_mmu_early_va_e[0]), .A1(byp_alu_rs1_data_e[0]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[0]) );
  HDMUX2D1 U657 ( .A0(exu_mmu_early_va_e[1]), .A1(byp_alu_rs1_data_e[1]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[1]) );
  HDMUX2D1 U646 ( .A0(exu_mmu_early_va_e[2]), .A1(byp_alu_rs1_data_e[2]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[2]) );
  HDMUX2D1 U635 ( .A0(exu_lsu_early_va_e[3]), .A1(byp_alu_rs1_data_e[3]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[3]) );
  HDMUX2D1 U627 ( .A0(exu_lsu_early_va_e[4]), .A1(byp_alu_rs1_data_e[4]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[4]) );
  HDMUX2D1 U626 ( .A0(exu_lsu_early_va_e[5]), .A1(byp_alu_rs1_data_e[5]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[5]) );
  HDMUX2D1 U625 ( .A0(exu_lsu_early_va_e[6]), .A1(byp_alu_rs1_data_e[6]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[6]) );
  HDMUX2D1 U624 ( .A0(exu_lsu_early_va_e[7]), .A1(byp_alu_rs1_data_e[7]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[7]) );
  HDMUX2D1 U623 ( .A0(exu_lsu_early_va_e[8]), .A1(byp_alu_rs1_data_e[8]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[8]) );
  HDMUX2D1 U622 ( .A0(exu_lsu_early_va_e[9]), .A1(byp_alu_rs1_data_e[9]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[9]) );
  HDMUX2D1 U667 ( .A0(exu_lsu_early_va_e[10]), .A1(byp_alu_rs1_data_e[10]), 
        .SL(ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[10]) );
  HDMUX2D1 U666 ( .A0(exu_ifu_brpc_e[11]), .A1(byp_alu_rs1_data_e[11]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[11]) );
  HDMUX2D1 U665 ( .A0(exu_ifu_brpc_e[12]), .A1(byp_alu_rs1_data_e[12]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[12]) );
  HDMUX2D1 U664 ( .A0(exu_ifu_brpc_e[13]), .A1(byp_alu_rs1_data_e[13]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[13]) );
  HDMUX2D1 U663 ( .A0(exu_ifu_brpc_e[14]), .A1(byp_alu_rs1_data_e[14]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[14]) );
  HDMUX2D1 U662 ( .A0(exu_ifu_brpc_e[15]), .A1(byp_alu_rs1_data_e[15]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[15]) );
  HDMUX2D1 U661 ( .A0(exu_ifu_brpc_e[16]), .A1(byp_alu_rs1_data_e[16]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[16]) );
  HDMUX2D1 U660 ( .A0(exu_ifu_brpc_e[17]), .A1(byp_alu_rs1_data_e[17]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[17]) );
  HDMUX2D1 U659 ( .A0(exu_ifu_brpc_e[18]), .A1(byp_alu_rs1_data_e[18]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[18]) );
  HDMUX2D1 U658 ( .A0(exu_ifu_brpc_e[19]), .A1(byp_alu_rs1_data_e[19]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[19]) );
  HDMUX2D1 U656 ( .A0(exu_ifu_brpc_e[20]), .A1(byp_alu_rs1_data_e[20]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[20]) );
  HDMUX2D1 U655 ( .A0(exu_ifu_brpc_e[21]), .A1(byp_alu_rs1_data_e[21]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[21]) );
  HDMUX2D1 U654 ( .A0(exu_ifu_brpc_e[22]), .A1(byp_alu_rs1_data_e[22]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[22]) );
  HDMUX2D1 U653 ( .A0(exu_ifu_brpc_e[23]), .A1(byp_alu_rs1_data_e[23]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[23]) );
  HDMUX2D1 U652 ( .A0(exu_ifu_brpc_e[24]), .A1(byp_alu_rs1_data_e[24]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[24]) );
  HDMUX2D1 U651 ( .A0(exu_ifu_brpc_e[25]), .A1(byp_alu_rs1_data_e[25]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[25]) );
  HDMUX2D1 U650 ( .A0(exu_ifu_brpc_e[26]), .A1(byp_alu_rs1_data_e[26]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[26]) );
  HDMUX2D1 U649 ( .A0(exu_ifu_brpc_e[27]), .A1(byp_alu_rs1_data_e[27]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[27]) );
  HDMUX2D1 U648 ( .A0(exu_ifu_brpc_e[28]), .A1(byp_alu_rs1_data_e[28]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[28]) );
  HDMUX2D1 U647 ( .A0(exu_ifu_brpc_e[29]), .A1(byp_alu_rs1_data_e[29]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[29]) );
  HDMUX2D1 U645 ( .A0(exu_ifu_brpc_e[30]), .A1(byp_alu_rs1_data_e[30]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[30]) );
  HDMUX2D1 U644 ( .A0(exu_ifu_brpc_e_31_), .A1(byp_alu_rs1_data_e[31]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[31]) );
  HDMUX2D1 U643 ( .A0(exu_ifu_brpc_e[32]), .A1(byp_alu_rs1_data_e[32]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[32]) );
  HDAOI22D1 U867 ( .A1(shft_alu_shift_out_e[63]), .A2(n947), .B1(
        alu_ecl_adder_out_63_e), .B2(n30), .Z(n448) );
  HDNAN2D1 U131 ( .A1(byp_alu_rs3_data_e[63]), .A2(n939), .Z(n449) );
  HDOAI211D1 U866 ( .A1(n346), .A2(ecl_alu_out_sel_logic_e_l), .B(n448), .C(
        n449), .Z(alu_byp_rd_data_e[63]) );
  HDAOI22D1 U875 ( .A1(shft_alu_shift_out_e[61]), .A2(n947), .B1(adder_out[61]), .B2(n30), .Z(n462) );
  HDNAN2D1 U143 ( .A1(byp_alu_rs3_data_e[61]), .A2(n939), .Z(n463) );
  HDOAI211D1 U874 ( .A1(n364), .A2(ecl_alu_out_sel_logic_e_l), .B(n462), .C(
        n463), .Z(alu_byp_rd_data_e[61]) );
  HDAOI22D1 U879 ( .A1(shft_alu_shift_out_e[60]), .A2(n947), .B1(adder_out[60]), .B2(n30), .Z(n469) );
  HDNAN2D1 U149 ( .A1(byp_alu_rs3_data_e[60]), .A2(n939), .Z(n470) );
  HDOAI211D1 U878 ( .A1(n363), .A2(ecl_alu_out_sel_logic_e_l), .B(n469), .C(
        n470), .Z(alu_byp_rd_data_e[60]) );
  HDAOI22D1 U887 ( .A1(shft_alu_shift_out_e[59]), .A2(n947), .B1(adder_out[59]), .B2(n30), .Z(n483) );
  HDNAN2D1 U161 ( .A1(byp_alu_rs3_data_e[59]), .A2(n939), .Z(n484) );
  HDOAI211D1 U886 ( .A1(n362), .A2(ecl_alu_out_sel_logic_e_l), .B(n483), .C(
        n484), .Z(alu_byp_rd_data_e[59]) );
  HDAOI22D1 U891 ( .A1(shft_alu_shift_out_e[58]), .A2(n947), .B1(adder_out[58]), .B2(n30), .Z(n490) );
  HDNAN2D1 U167 ( .A1(byp_alu_rs3_data_e[58]), .A2(n939), .Z(n491) );
  HDOAI211D1 U890 ( .A1(n361), .A2(ecl_alu_out_sel_logic_e_l), .B(n490), .C(
        n491), .Z(alu_byp_rd_data_e[58]) );
  HDAOI22D1 U895 ( .A1(shft_alu_shift_out_e[57]), .A2(n947), .B1(adder_out[57]), .B2(n30), .Z(n497) );
  HDNAN2D1 U173 ( .A1(byp_alu_rs3_data_e[57]), .A2(n939), .Z(n498) );
  HDOAI211D1 U894 ( .A1(n360), .A2(ecl_alu_out_sel_logic_e_l), .B(n497), .C(
        n498), .Z(alu_byp_rd_data_e[57]) );
  HDAOI22D1 U899 ( .A1(shft_alu_shift_out_e[56]), .A2(n947), .B1(adder_out[56]), .B2(n30), .Z(n504) );
  HDNAN2D1 U179 ( .A1(byp_alu_rs3_data_e[56]), .A2(n939), .Z(n505) );
  HDOAI211D1 U898 ( .A1(n359), .A2(ecl_alu_out_sel_logic_e_l), .B(n504), .C(
        n505), .Z(alu_byp_rd_data_e[56]) );
  HDAOI22D1 U903 ( .A1(shft_alu_shift_out_e[55]), .A2(n947), .B1(adder_out[55]), .B2(n30), .Z(n511) );
  HDNAN2D1 U185 ( .A1(byp_alu_rs3_data_e[55]), .A2(n939), .Z(n512) );
  HDOAI211D1 U902 ( .A1(n358), .A2(ecl_alu_out_sel_logic_e_l), .B(n511), .C(
        n512), .Z(alu_byp_rd_data_e[55]) );
  HDAOI22D1 U907 ( .A1(shft_alu_shift_out_e[54]), .A2(n946), .B1(adder_out[54]), .B2(n30), .Z(n518) );
  HDNAN2D1 U191 ( .A1(byp_alu_rs3_data_e[54]), .A2(n939), .Z(n519) );
  HDOAI211D1 U906 ( .A1(n373), .A2(ecl_alu_out_sel_logic_e_l), .B(n518), .C(
        n519), .Z(alu_byp_rd_data_e[54]) );
  HDAOI22D1 U911 ( .A1(shft_alu_shift_out_e[53]), .A2(n946), .B1(adder_out[53]), .B2(n30), .Z(n525) );
  HDNAN2D1 U197 ( .A1(byp_alu_rs3_data_e[53]), .A2(n939), .Z(n526) );
  HDOAI211D1 U910 ( .A1(n372), .A2(ecl_alu_out_sel_logic_e_l), .B(n525), .C(
        n526), .Z(alu_byp_rd_data_e[53]) );
  HDAOI22D1 U915 ( .A1(shft_alu_shift_out_e[52]), .A2(n946), .B1(adder_out[52]), .B2(n30), .Z(n532) );
  HDNAN2D1 U203 ( .A1(byp_alu_rs3_data_e[52]), .A2(n939), .Z(n533) );
  HDOAI211D1 U914 ( .A1(n371), .A2(ecl_alu_out_sel_logic_e_l), .B(n532), .C(
        n533), .Z(alu_byp_rd_data_e[52]) );
  HDAOI22D1 U919 ( .A1(shft_alu_shift_out_e[51]), .A2(n946), .B1(adder_out[51]), .B2(n30), .Z(n539) );
  HDNAN2D1 U209 ( .A1(byp_alu_rs3_data_e[51]), .A2(n939), .Z(n540) );
  HDOAI211D1 U918 ( .A1(n370), .A2(ecl_alu_out_sel_logic_e_l), .B(n539), .C(
        n540), .Z(alu_byp_rd_data_e[51]) );
  HDAOI22D1 U923 ( .A1(shft_alu_shift_out_e[50]), .A2(n946), .B1(adder_out[50]), .B2(n952), .Z(n546) );
  HDNAN2D1 U215 ( .A1(byp_alu_rs3_data_e[50]), .A2(n939), .Z(n547) );
  HDOAI211D1 U922 ( .A1(n369), .A2(ecl_alu_out_sel_logic_e_l), .B(n546), .C(
        n547), .Z(alu_byp_rd_data_e[50]) );
  HDAOI22D1 U931 ( .A1(shft_alu_shift_out_e[49]), .A2(n946), .B1(adder_out[49]), .B2(n952), .Z(n560) );
  HDNAN2D1 U227 ( .A1(byp_alu_rs3_data_e[49]), .A2(n939), .Z(n561) );
  HDOAI211D1 U930 ( .A1(n368), .A2(ecl_alu_out_sel_logic_e_l), .B(n560), .C(
        n561), .Z(alu_byp_rd_data_e[49]) );
  HDAOI22D1 U935 ( .A1(shft_alu_shift_out_e[48]), .A2(n946), .B1(adder_out[48]), .B2(n952), .Z(n567) );
  HDNAN2D1 U233 ( .A1(byp_alu_rs3_data_e[48]), .A2(n939), .Z(n568) );
  HDOAI211D1 U934 ( .A1(n367), .A2(ecl_alu_out_sel_logic_e_l), .B(n567), .C(
        n568), .Z(alu_byp_rd_data_e[48]) );
  HDAOI22D1 U939 ( .A1(byp_alu_rs3_data_e[47]), .A2(n417), .B1(
        exu_ifu_brpc_e[47]), .B2(n952), .Z(n574) );
  HDNAN2D1 U239 ( .A1(shft_alu_shift_out_e[47]), .A2(n942), .Z(n575) );
  HDOAI211D1 U938 ( .A1(n366), .A2(ecl_alu_out_sel_logic_e_l), .B(n574), .C(
        n575), .Z(alu_byp_rd_data_e[47]) );
  HDAOI22D1 U943 ( .A1(byp_alu_rs3_data_e[46]), .A2(n417), .B1(
        exu_ifu_brpc_e[46]), .B2(n952), .Z(n581) );
  HDNAN2D1 U245 ( .A1(shft_alu_shift_out_e[46]), .A2(n945), .Z(n582) );
  HDOAI211D1 U942 ( .A1(n345), .A2(ecl_alu_out_sel_logic_e_l), .B(n581), .C(
        n582), .Z(alu_byp_rd_data_e[46]) );
  HDAOI22D1 U947 ( .A1(byp_alu_rs3_data_e[45]), .A2(n417), .B1(
        exu_ifu_brpc_e[45]), .B2(n952), .Z(n588) );
  HDNAN2D1 U251 ( .A1(shft_alu_shift_out_e[45]), .A2(n944), .Z(n589) );
  HDOAI211D1 U946 ( .A1(n344), .A2(ecl_alu_out_sel_logic_e_l), .B(n588), .C(
        n589), .Z(alu_byp_rd_data_e[45]) );
  HDAOI22D1 U951 ( .A1(byp_alu_rs3_data_e[44]), .A2(n417), .B1(
        exu_ifu_brpc_e[44]), .B2(n952), .Z(n595) );
  HDNAN2D1 U257 ( .A1(shft_alu_shift_out_e[44]), .A2(n943), .Z(n596) );
  HDOAI211D1 U950 ( .A1(n343), .A2(ecl_alu_out_sel_logic_e_l), .B(n595), .C(
        n596), .Z(alu_byp_rd_data_e[44]) );
  HDAOI22D1 U955 ( .A1(byp_alu_rs3_data_e[43]), .A2(n417), .B1(
        exu_ifu_brpc_e[43]), .B2(n951), .Z(n602) );
  HDNAN2D1 U263 ( .A1(shft_alu_shift_out_e[43]), .A2(n942), .Z(n603) );
  HDOAI211D1 U954 ( .A1(n342), .A2(ecl_alu_out_sel_logic_e_l), .B(n602), .C(
        n603), .Z(alu_byp_rd_data_e[43]) );
  HDAOI22D1 U959 ( .A1(byp_alu_rs3_data_e[42]), .A2(n417), .B1(
        exu_ifu_brpc_e[42]), .B2(n951), .Z(n609) );
  HDNAN2D1 U269 ( .A1(shft_alu_shift_out_e[42]), .A2(n947), .Z(n610) );
  HDOAI211D1 U958 ( .A1(n341), .A2(ecl_alu_out_sel_logic_e_l), .B(n609), .C(
        n610), .Z(alu_byp_rd_data_e[42]) );
  HDAOI22D1 U963 ( .A1(byp_alu_rs3_data_e[41]), .A2(n417), .B1(
        exu_ifu_brpc_e[41]), .B2(n951), .Z(n616) );
  HDNAN2D1 U275 ( .A1(shft_alu_shift_out_e[41]), .A2(n945), .Z(n617) );
  HDOAI211D1 U962 ( .A1(n340), .A2(ecl_alu_out_sel_logic_e_l), .B(n616), .C(
        n617), .Z(alu_byp_rd_data_e[41]) );
  HDAOI22D1 U967 ( .A1(byp_alu_rs3_data_e[40]), .A2(n417), .B1(
        exu_ifu_brpc_e[40]), .B2(n951), .Z(n623) );
  HDNAN2D1 U281 ( .A1(shft_alu_shift_out_e[40]), .A2(n945), .Z(n624) );
  HDOAI211D1 U966 ( .A1(n339), .A2(ecl_alu_out_sel_logic_e_l), .B(n623), .C(
        n624), .Z(alu_byp_rd_data_e[40]) );
  HDAOI22D1 U975 ( .A1(byp_alu_rs3_data_e[39]), .A2(n417), .B1(
        exu_ifu_brpc_e[39]), .B2(n951), .Z(n637) );
  HDNAN2D1 U293 ( .A1(shft_alu_shift_out_e[39]), .A2(n945), .Z(n638) );
  HDOAI211D1 U974 ( .A1(n338), .A2(ecl_alu_out_sel_logic_e_l), .B(n637), .C(
        n638), .Z(alu_byp_rd_data_e[39]) );
  HDAOI22D1 U979 ( .A1(byp_alu_rs3_data_e[38]), .A2(n417), .B1(
        exu_ifu_brpc_e[38]), .B2(n951), .Z(n644) );
  HDNAN2D1 U299 ( .A1(shft_alu_shift_out_e[38]), .A2(n945), .Z(n645) );
  HDOAI211D1 U978 ( .A1(n353), .A2(ecl_alu_out_sel_logic_e_l), .B(n644), .C(
        n645), .Z(alu_byp_rd_data_e[38]) );
  HDAOI22D1 U983 ( .A1(byp_alu_rs3_data_e[37]), .A2(n417), .B1(
        exu_ifu_brpc_e[37]), .B2(n951), .Z(n651) );
  HDNAN2D1 U305 ( .A1(shft_alu_shift_out_e[37]), .A2(n945), .Z(n652) );
  HDOAI211D1 U982 ( .A1(n352), .A2(ecl_alu_out_sel_logic_e_l), .B(n651), .C(
        n652), .Z(alu_byp_rd_data_e[37]) );
  HDAOI22D1 U987 ( .A1(byp_alu_rs3_data_e[36]), .A2(n417), .B1(
        exu_ifu_brpc_e[36]), .B2(n950), .Z(n658) );
  HDNAN2D1 U311 ( .A1(shft_alu_shift_out_e[36]), .A2(n945), .Z(n659) );
  HDOAI211D1 U986 ( .A1(n351), .A2(ecl_alu_out_sel_logic_e_l), .B(n658), .C(
        n659), .Z(alu_byp_rd_data_e[36]) );
  HDAOI22D1 U991 ( .A1(byp_alu_rs3_data_e[35]), .A2(n417), .B1(
        exu_ifu_brpc_e[35]), .B2(n950), .Z(n665) );
  HDNAN2D1 U317 ( .A1(shft_alu_shift_out_e[35]), .A2(n945), .Z(n666) );
  HDOAI211D1 U990 ( .A1(n350), .A2(ecl_alu_out_sel_logic_e_l), .B(n665), .C(
        n666), .Z(alu_byp_rd_data_e[35]) );
  HDAOI22D1 U995 ( .A1(byp_alu_rs3_data_e[34]), .A2(n417), .B1(
        exu_ifu_brpc_e[34]), .B2(n950), .Z(n672) );
  HDNAN2D1 U323 ( .A1(shft_alu_shift_out_e[34]), .A2(n945), .Z(n673) );
  HDOAI211D1 U994 ( .A1(n349), .A2(ecl_alu_out_sel_logic_e_l), .B(n672), .C(
        n673), .Z(alu_byp_rd_data_e[34]) );
  HDAOI22D1 U999 ( .A1(byp_alu_rs3_data_e[33]), .A2(n417), .B1(
        exu_ifu_brpc_e[33]), .B2(n950), .Z(n679) );
  HDNAN2D1 U329 ( .A1(shft_alu_shift_out_e[33]), .A2(n944), .Z(n680) );
  HDOAI211D1 U998 ( .A1(n348), .A2(ecl_alu_out_sel_logic_e_l), .B(n679), .C(
        n680), .Z(alu_byp_rd_data_e[33]) );
  HDAOI22D1 U1003 ( .A1(byp_alu_rs3_data_e[32]), .A2(n417), .B1(
        exu_ifu_brpc_e[32]), .B2(n950), .Z(n686) );
  HDNAN2D1 U335 ( .A1(shft_alu_shift_out_e[32]), .A2(n944), .Z(n687) );
  HDOAI211D1 U1002 ( .A1(n347), .A2(ecl_alu_out_sel_logic_e_l), .B(n686), .C(
        n687), .Z(alu_byp_rd_data_e[32]) );
  HDAOI22D1 U1008 ( .A1(byp_alu_rs3_data_e[31]), .A2(n417), .B1(
        exu_ifu_brpc_e_31_), .B2(n950), .Z(n693) );
  HDNAN2D1 U341 ( .A1(shft_alu_shift_out_e[31]), .A2(n944), .Z(n694) );
  HDOAI211D1 U1007 ( .A1(n173), .A2(ecl_alu_out_sel_logic_e_l), .B(n693), .C(
        n694), .Z(alu_byp_rd_data_e[31]) );
  HDAOI22D1 U1013 ( .A1(byp_alu_rs3_data_e[30]), .A2(n417), .B1(
        exu_ifu_brpc_e[30]), .B2(n950), .Z(n700) );
  HDNAN2D1 U347 ( .A1(shft_alu_shift_out_e[30]), .A2(n944), .Z(n701) );
  HDOAI211D1 U1012 ( .A1(n192), .A2(ecl_alu_out_sel_logic_e_l), .B(n700), .C(
        n701), .Z(alu_byp_rd_data_e[30]) );
  HDAOI22D1 U1021 ( .A1(byp_alu_rs3_data_e[29]), .A2(n417), .B1(
        exu_ifu_brpc_e[29]), .B2(n949), .Z(n714) );
  HDNAN2D1 U359 ( .A1(shft_alu_shift_out_e[29]), .A2(n944), .Z(n715) );
  HDOAI211D1 U1020 ( .A1(n191), .A2(ecl_alu_out_sel_logic_e_l), .B(n714), .C(
        n715), .Z(alu_byp_rd_data_e[29]) );
  HDAOI22D1 U1025 ( .A1(byp_alu_rs3_data_e[28]), .A2(n939), .B1(
        exu_ifu_brpc_e[28]), .B2(n949), .Z(n721) );
  HDNAN2D1 U365 ( .A1(shft_alu_shift_out_e[28]), .A2(n944), .Z(n722) );
  HDOAI211D1 U1024 ( .A1(n190), .A2(ecl_alu_out_sel_logic_e_l), .B(n721), .C(
        n722), .Z(alu_byp_rd_data_e[28]) );
  HDAOI22D1 U1029 ( .A1(byp_alu_rs3_data_e[27]), .A2(n939), .B1(
        exu_ifu_brpc_e[27]), .B2(n949), .Z(n728) );
  HDNAN2D1 U371 ( .A1(shft_alu_shift_out_e[27]), .A2(n944), .Z(n729) );
  HDOAI211D1 U1028 ( .A1(n189), .A2(ecl_alu_out_sel_logic_e_l), .B(n728), .C(
        n729), .Z(alu_byp_rd_data_e[27]) );
  HDAOI22D1 U1033 ( .A1(byp_alu_rs3_data_e[26]), .A2(n939), .B1(
        exu_ifu_brpc_e[26]), .B2(n949), .Z(n735) );
  HDNAN2D1 U377 ( .A1(shft_alu_shift_out_e[26]), .A2(n944), .Z(n736) );
  HDOAI211D1 U1032 ( .A1(n188), .A2(ecl_alu_out_sel_logic_e_l), .B(n735), .C(
        n736), .Z(alu_byp_rd_data_e[26]) );
  HDAOI22D1 U1037 ( .A1(byp_alu_rs3_data_e[25]), .A2(n939), .B1(
        exu_ifu_brpc_e[25]), .B2(n949), .Z(n742) );
  HDNAN2D1 U383 ( .A1(shft_alu_shift_out_e[25]), .A2(n943), .Z(n743) );
  HDOAI211D1 U1036 ( .A1(n187), .A2(ecl_alu_out_sel_logic_e_l), .B(n742), .C(
        n743), .Z(alu_byp_rd_data_e[25]) );
  HDAOI22D1 U1041 ( .A1(byp_alu_rs3_data_e[24]), .A2(n939), .B1(
        exu_ifu_brpc_e[24]), .B2(n949), .Z(n749) );
  HDNAN2D1 U389 ( .A1(shft_alu_shift_out_e[24]), .A2(n943), .Z(n750) );
  HDOAI211D1 U1040 ( .A1(n186), .A2(ecl_alu_out_sel_logic_e_l), .B(n749), .C(
        n750), .Z(alu_byp_rd_data_e[24]) );
  HDAOI22D1 U1045 ( .A1(byp_alu_rs3_data_e[23]), .A2(n939), .B1(
        exu_ifu_brpc_e[23]), .B2(n949), .Z(n756) );
  HDNAN2D1 U395 ( .A1(shft_alu_shift_out_e[23]), .A2(n943), .Z(n757) );
  HDOAI211D1 U1044 ( .A1(n185), .A2(ecl_alu_out_sel_logic_e_l), .B(n756), .C(
        n757), .Z(alu_byp_rd_data_e[23]) );
  HDAOI22D1 U1049 ( .A1(byp_alu_rs3_data_e[22]), .A2(n939), .B1(
        exu_ifu_brpc_e[22]), .B2(n949), .Z(n763) );
  HDNAN2D1 U401 ( .A1(shft_alu_shift_out_e[22]), .A2(n943), .Z(n764) );
  HDOAI211D1 U1048 ( .A1(n200), .A2(ecl_alu_out_sel_logic_e_l), .B(n763), .C(
        n764), .Z(alu_byp_rd_data_e[22]) );
  HDAOI22D1 U1053 ( .A1(byp_alu_rs3_data_e[21]), .A2(n417), .B1(
        exu_ifu_brpc_e[21]), .B2(n948), .Z(n770) );
  HDNAN2D1 U407 ( .A1(shft_alu_shift_out_e[21]), .A2(n943), .Z(n771) );
  HDOAI211D1 U1052 ( .A1(n199), .A2(ecl_alu_out_sel_logic_e_l), .B(n770), .C(
        n771), .Z(alu_byp_rd_data_e[21]) );
  HDAOI22D1 U1057 ( .A1(byp_alu_rs3_data_e[20]), .A2(n939), .B1(
        exu_ifu_brpc_e[20]), .B2(n948), .Z(n777) );
  HDNAN2D1 U413 ( .A1(shft_alu_shift_out_e[20]), .A2(n943), .Z(n778) );
  HDOAI211D1 U1056 ( .A1(n198), .A2(ecl_alu_out_sel_logic_e_l), .B(n777), .C(
        n778), .Z(alu_byp_rd_data_e[20]) );
  HDAOI22D1 U1065 ( .A1(byp_alu_rs3_data_e[19]), .A2(n417), .B1(
        exu_ifu_brpc_e[19]), .B2(n948), .Z(n791) );
  HDNAN2D1 U425 ( .A1(shft_alu_shift_out_e[19]), .A2(n943), .Z(n792) );
  HDOAI211D1 U1064 ( .A1(n197), .A2(ecl_alu_out_sel_logic_e_l), .B(n791), .C(
        n792), .Z(alu_byp_rd_data_e[19]) );
  HDAOI22D1 U1069 ( .A1(byp_alu_rs3_data_e[18]), .A2(n417), .B1(
        exu_ifu_brpc_e[18]), .B2(n948), .Z(n798) );
  HDNAN2D1 U431 ( .A1(shft_alu_shift_out_e[18]), .A2(n943), .Z(n799) );
  HDOAI211D1 U1068 ( .A1(n196), .A2(ecl_alu_out_sel_logic_e_l), .B(n798), .C(
        n799), .Z(alu_byp_rd_data_e[18]) );
  HDAOI22D1 U1073 ( .A1(byp_alu_rs3_data_e[17]), .A2(n417), .B1(
        exu_ifu_brpc_e[17]), .B2(n948), .Z(n805) );
  HDNAN2D1 U437 ( .A1(shft_alu_shift_out_e[17]), .A2(n942), .Z(n806) );
  HDOAI211D1 U1072 ( .A1(n195), .A2(ecl_alu_out_sel_logic_e_l), .B(n805), .C(
        n806), .Z(alu_byp_rd_data_e[17]) );
  HDAOI22D1 U1077 ( .A1(byp_alu_rs3_data_e[16]), .A2(n417), .B1(
        exu_ifu_brpc_e[16]), .B2(n948), .Z(n812) );
  HDNAN2D1 U443 ( .A1(shft_alu_shift_out_e[16]), .A2(n942), .Z(n813) );
  HDOAI211D1 U1076 ( .A1(n194), .A2(ecl_alu_out_sel_logic_e_l), .B(n812), .C(
        n813), .Z(alu_byp_rd_data_e[16]) );
  HDAOI22D1 U1081 ( .A1(byp_alu_rs3_data_e[15]), .A2(n417), .B1(
        exu_ifu_brpc_e[15]), .B2(n948), .Z(n819) );
  HDNAN2D1 U449 ( .A1(shft_alu_shift_out_e[15]), .A2(n942), .Z(n820) );
  HDOAI211D1 U1080 ( .A1(n193), .A2(ecl_alu_out_sel_logic_e_l), .B(n819), .C(
        n820), .Z(alu_byp_rd_data_e[15]) );
  HDAOI22D1 U1085 ( .A1(byp_alu_rs3_data_e[14]), .A2(n417), .B1(
        exu_ifu_brpc_e[14]), .B2(n951), .Z(n826) );
  HDNAN2D1 U455 ( .A1(shft_alu_shift_out_e[14]), .A2(n942), .Z(n827) );
  HDOAI211D1 U1084 ( .A1(n172), .A2(ecl_alu_out_sel_logic_e_l), .B(n826), .C(
        n827), .Z(alu_byp_rd_data_e[14]) );
  HDAOI22D1 U1089 ( .A1(byp_alu_rs3_data_e[13]), .A2(n417), .B1(
        exu_ifu_brpc_e[13]), .B2(n950), .Z(n833) );
  HDNAN2D1 U461 ( .A1(shft_alu_shift_out_e[13]), .A2(n942), .Z(n834) );
  HDOAI211D1 U1088 ( .A1(n171), .A2(ecl_alu_out_sel_logic_e_l), .B(n833), .C(
        n834), .Z(alu_byp_rd_data_e[13]) );
  HDAOI22D1 U1093 ( .A1(byp_alu_rs3_data_e[12]), .A2(n417), .B1(
        exu_ifu_brpc_e[12]), .B2(n952), .Z(n840) );
  HDNAN2D1 U467 ( .A1(shft_alu_shift_out_e[12]), .A2(n942), .Z(n841) );
  HDOAI211D1 U1092 ( .A1(n170), .A2(ecl_alu_out_sel_logic_e_l), .B(n840), .C(
        n841), .Z(alu_byp_rd_data_e[12]) );
  HDAOI22D1 U1097 ( .A1(byp_alu_rs3_data_e[11]), .A2(n417), .B1(
        exu_ifu_brpc_e[11]), .B2(n952), .Z(n847) );
  HDNAN2D1 U473 ( .A1(shft_alu_shift_out_e[11]), .A2(n942), .Z(n848) );
  HDOAI211D1 U1096 ( .A1(n169), .A2(ecl_alu_out_sel_logic_e_l), .B(n847), .C(
        n848), .Z(alu_byp_rd_data_e[11]) );
  HDAOI22D1 U1101 ( .A1(byp_alu_rs3_data_e[10]), .A2(n939), .B1(
        exu_lsu_early_va_e[10]), .B2(n949), .Z(n854) );
  HDNAN2D1 U479 ( .A1(shft_alu_shift_out_e[10]), .A2(n942), .Z(n855) );
  HDOAI211D1 U1100 ( .A1(n168), .A2(ecl_alu_out_sel_logic_e_l), .B(n854), .C(
        n855), .Z(alu_byp_rd_data_e[10]) );
  HDAOI22D1 U851 ( .A1(byp_alu_rs3_data_e[9]), .A2(n417), .B1(
        exu_lsu_early_va_e[9]), .B2(n30), .Z(n414) );
  HDNAN2D1 U107 ( .A1(shft_alu_shift_out_e[9]), .A2(n946), .Z(n415) );
  HDOAI211D1 U850 ( .A1(n167), .A2(ecl_alu_out_sel_logic_e_l), .B(n414), .C(
        n415), .Z(alu_byp_rd_data_e[9]) );
  HDAOI22D1 U855 ( .A1(byp_alu_rs3_data_e[8]), .A2(n417), .B1(
        exu_lsu_early_va_e[8]), .B2(n30), .Z(n427) );
  HDNAN2D1 U113 ( .A1(shft_alu_shift_out_e[8]), .A2(n946), .Z(n428) );
  HDOAI211D1 U854 ( .A1(n166), .A2(ecl_alu_out_sel_logic_e_l), .B(n427), .C(
        n428), .Z(alu_byp_rd_data_e[8]) );
  HDAOI22D1 U859 ( .A1(byp_alu_rs3_data_e[7]), .A2(n417), .B1(
        exu_lsu_early_va_e[7]), .B2(n30), .Z(n434) );
  HDNAN2D1 U119 ( .A1(shft_alu_shift_out_e[7]), .A2(n946), .Z(n435) );
  HDOAI211D1 U858 ( .A1(n165), .A2(ecl_alu_out_sel_logic_e_l), .B(n434), .C(
        n435), .Z(alu_byp_rd_data_e[7]) );
  HDAOI22D1 U863 ( .A1(byp_alu_rs3_data_e[6]), .A2(n417), .B1(
        exu_lsu_early_va_e[6]), .B2(n30), .Z(n441) );
  HDNAN2D1 U125 ( .A1(shft_alu_shift_out_e[6]), .A2(n945), .Z(n442) );
  HDOAI211D1 U862 ( .A1(n180), .A2(ecl_alu_out_sel_logic_e_l), .B(n441), .C(
        n442), .Z(alu_byp_rd_data_e[6]) );
  HDAOI22D1 U883 ( .A1(byp_alu_rs3_data_e[5]), .A2(n417), .B1(
        exu_lsu_early_va_e[5]), .B2(n30), .Z(n476) );
  HDNAN2D1 U155 ( .A1(shft_alu_shift_out_e[5]), .A2(n944), .Z(n477) );
  HDOAI211D1 U882 ( .A1(n179), .A2(ecl_alu_out_sel_logic_e_l), .B(n476), .C(
        n477), .Z(alu_byp_rd_data_e[5]) );
  HDAOI22D1 U927 ( .A1(byp_alu_rs3_data_e[4]), .A2(n417), .B1(
        exu_lsu_early_va_e[4]), .B2(n952), .Z(n553) );
  HDNAN2D1 U221 ( .A1(shft_alu_shift_out_e[4]), .A2(n943), .Z(n554) );
  HDOAI211D1 U926 ( .A1(n178), .A2(ecl_alu_out_sel_logic_e_l), .B(n553), .C(
        n554), .Z(alu_byp_rd_data_e[4]) );
  HDAOI22D1 U971 ( .A1(byp_alu_rs3_data_e[3]), .A2(n417), .B1(
        exu_lsu_early_va_e[3]), .B2(n951), .Z(n630) );
  HDNAN2D1 U287 ( .A1(shft_alu_shift_out_e[3]), .A2(n945), .Z(n631) );
  HDOAI211D1 U970 ( .A1(n177), .A2(ecl_alu_out_sel_logic_e_l), .B(n630), .C(
        n631), .Z(alu_byp_rd_data_e[3]) );
  HDAOI22D1 U1017 ( .A1(byp_alu_rs3_data_e[2]), .A2(n417), .B1(
        exu_mmu_early_va_e[2]), .B2(n950), .Z(n707) );
  HDNAN2D1 U353 ( .A1(shft_alu_shift_out_e[2]), .A2(n944), .Z(n708) );
  HDOAI211D1 U1016 ( .A1(n176), .A2(ecl_alu_out_sel_logic_e_l), .B(n707), .C(
        n708), .Z(alu_byp_rd_data_e[2]) );
  HDAOI22D1 U1061 ( .A1(byp_alu_rs3_data_e[1]), .A2(n417), .B1(
        exu_mmu_early_va_e[1]), .B2(n948), .Z(n784) );
  HDNAN2D1 U419 ( .A1(shft_alu_shift_out_e[1]), .A2(n943), .Z(n785) );
  HDOAI211D1 U1060 ( .A1(n175), .A2(ecl_alu_out_sel_logic_e_l), .B(n784), .C(
        n785), .Z(alu_byp_rd_data_e[1]) );
  HDAOI22D1 U1105 ( .A1(byp_alu_rs3_data_e[0]), .A2(n939), .B1(
        exu_mmu_early_va_e[0]), .B2(n948), .Z(n861) );
  HDNAN2D1 U485 ( .A1(shft_alu_shift_out_e[0]), .A2(n942), .Z(n862) );
  HDOAI211D1 U1104 ( .A1(n174), .A2(ecl_alu_out_sel_logic_e_l), .B(n861), .C(
        n862), .Z(alu_byp_rd_data_e[0]) );
  HDMUX2D1 U642 ( .A0(exu_ifu_brpc_e[33]), .A1(byp_alu_rs1_data_e[33]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[33]) );
  HDMUX2D1 U628 ( .A0(exu_ifu_brpc_e[46]), .A1(byp_alu_rs1_data_e[46]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[46]) );
  HDMUX2D1 U629 ( .A0(exu_ifu_brpc_e[45]), .A1(byp_alu_rs1_data_e[45]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[45]) );
  HDMUX2D1 U630 ( .A0(exu_ifu_brpc_e[44]), .A1(byp_alu_rs1_data_e[44]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[44]) );
  HDMUX2D1 U631 ( .A0(exu_ifu_brpc_e[43]), .A1(byp_alu_rs1_data_e[43]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[43]) );
  HDMUX2D1 U632 ( .A0(exu_ifu_brpc_e[42]), .A1(byp_alu_rs1_data_e[42]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[42]) );
  HDMUX2D1 U633 ( .A0(exu_ifu_brpc_e[41]), .A1(byp_alu_rs1_data_e[41]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[41]) );
  HDMUX2D1 U634 ( .A0(exu_ifu_brpc_e[40]), .A1(byp_alu_rs1_data_e[40]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[40]) );
  HDMUX2D1 U636 ( .A0(exu_ifu_brpc_e[39]), .A1(byp_alu_rs1_data_e[39]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[39]) );
  HDMUX2D1 U637 ( .A0(exu_ifu_brpc_e[38]), .A1(byp_alu_rs1_data_e[38]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[38]) );
  HDMUX2D1 U638 ( .A0(exu_ifu_brpc_e[37]), .A1(byp_alu_rs1_data_e[37]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[37]) );
  HDMUX2D1 U639 ( .A0(exu_ifu_brpc_e[36]), .A1(byp_alu_rs1_data_e[36]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[36]) );
  HDMUX2D1 U640 ( .A0(exu_ifu_brpc_e[35]), .A1(byp_alu_rs1_data_e[35]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[35]) );
  HDMUX2D1 U641 ( .A0(exu_ifu_brpc_e[34]), .A1(byp_alu_rs1_data_e[34]), .SL(
        ifu_lsu_casa_e), .Z(exu_lsu_ldst_va_e[34]) );
  HDAOI22D1 U871 ( .A1(shft_alu_shift_out_e[62]), .A2(n947), .B1(adder_out[62]), .B2(n30), .Z(n455) );
  HDNAN2D1 U137 ( .A1(byp_alu_rs3_data_e[62]), .A2(n939), .Z(n456) );
  HDOAI211D1 U870 ( .A1(n365), .A2(ecl_alu_out_sel_logic_e_l), .B(n455), .C(
        n456), .Z(alu_byp_rd_data_e[62]) );
  HDMUXB2DL U604 ( .A0(byp_alu_rs2_data_e_l[40]), .A1(n921), .SL(
        addsub_subtract_e[40]), .Z(addsub_rs2_data_40_) );
  HDMUXB2DL U608 ( .A0(byp_alu_rs2_data_e_l[38]), .A1(n923), .SL(
        addsub_subtract_e[38]), .Z(addsub_rs2_data_38_) );
  HDMUXB2DL U616 ( .A0(byp_alu_rs2_data_e_l[34]), .A1(n927), .SL(
        addsub_subtract_e[34]), .Z(addsub_rs2_data_34_) );
  HDMUXB2DL U618 ( .A0(byp_alu_rs2_data_e_l[33]), .A1(n928), .SL(
        addsub_subtract_e[33]), .Z(addsub_rs2_data_33_) );
  HDMUXB2DL U620 ( .A0(byp_alu_rs2_data_e_l[32]), .A1(n929), .SL(
        addsub_subtract_e[32]), .Z(addsub_rs2_data_32_) );
  HDMUXB2DL U522 ( .A0(byp_alu_rs2_data_e_l[25]), .A1(n880), .SL(
        addsub_subtract_e[25]), .Z(addsub_rs2_data_25) );
  HDMUXB2DL U524 ( .A0(byp_alu_rs2_data_e_l[24]), .A1(n881), .SL(
        addsub_subtract_e[24]), .Z(addsub_rs2_data_24) );
  HDMUXB2DL U526 ( .A0(byp_alu_rs2_data_e_l[23]), .A1(n882), .SL(
        addsub_subtract_e[23]), .Z(addsub_rs2_data_23) );
  HDMUXB2DL U528 ( .A0(byp_alu_rs2_data_e_l[22]), .A1(n883), .SL(
        addsub_subtract_e[22]), .Z(addsub_rs2_data_22) );
  HDMUXB2DL U530 ( .A0(byp_alu_rs2_data_e_l[21]), .A1(n884), .SL(
        addsub_subtract_e[21]), .Z(addsub_rs2_data_21) );
  HDMUXB2DL U532 ( .A0(byp_alu_rs2_data_e_l[20]), .A1(n885), .SL(
        addsub_subtract_e[20]), .Z(addsub_rs2_data_20) );
  HDMUXB2DL U550 ( .A0(byp_alu_rs2_data_e_l[12]), .A1(n894), .SL(
        addsub_subtract_e[12]), .Z(addsub_rs2_data_12) );
  HDMUXB2DL U552 ( .A0(byp_alu_rs2_data_e_l[11]), .A1(n895), .SL(
        addsub_subtract_e[11]), .Z(addsub_rs2_data_11) );
  HDMUXB2DL U554 ( .A0(byp_alu_rs2_data_e_l[10]), .A1(n896), .SL(
        addsub_subtract_e[10]), .Z(addsub_rs2_data_10) );
  HDMUXB2DL U508 ( .A0(byp_alu_rs2_data_e_l[4]), .A1(n873), .SL(
        addsub_subtract_e[4]), .Z(addsub_rs2_data_4) );
  HDMUXB2DL U512 ( .A0(byp_alu_rs2_data_e_l[3]), .A1(n875), .SL(
        addsub_subtract_e[3]), .Z(addsub_rs2_data_3) );
  HDNOR2D1 U94 ( .A1(n403), .A2(exu_lsu_ldst_va_e[47]), .Z(n411) );
  HDAOI211D1 U847 ( .A1(n403), .A2(exu_lsu_ldst_va_e[47]), .B(n410), .C(n411), 
        .Z(n409) );
  HDNAN4D1 U760 ( .A1(n197), .A2(n198), .A3(n199), .A4(n200), .Z(n181) );
  HDNAN4D1 U759 ( .A1(n193), .A2(n194), .A3(n195), .A4(n196), .Z(n182) );
  HDNAN4D1 U758 ( .A1(n189), .A2(n190), .A3(n191), .A4(n192), .Z(n183) );
  HDNAN4D1 U757 ( .A1(n185), .A2(n186), .A3(n187), .A4(n188), .Z(n184) );
  HDNAN4D1 U755 ( .A1(n177), .A2(n178), .A3(n179), .A4(n180), .Z(n161) );
  HDNAN4D1 U754 ( .A1(n173), .A2(n174), .A3(n175), .A4(n176), .Z(n162) );
  HDNAN4D1 U753 ( .A1(n169), .A2(n170), .A3(n171), .A4(n172), .Z(n163) );
  HDNAN4D1 U752 ( .A1(n165), .A2(n166), .A3(n167), .A4(n168), .Z(n164) );
  HDAO32DL U3 ( .A1(n28), .A2(n29), .A3(ecl_alu_out_sel_sum_e_l), .B1(n950), 
        .B2(n31), .Z(alu_ecl_zlow_e) );
  HDNAN2M1D1 U1005 ( .A1(ecl_alu_sethi_inst_e), .A2(ecl_alu_log_sel_move_e), 
        .Z(n450) );
  HDNAN4D1 U835 ( .A1(n370), .A2(n371), .A3(n372), .A4(n373), .Z(n354) );
  HDNAN4D1 U834 ( .A1(n366), .A2(n367), .A3(n368), .A4(n369), .Z(n355) );
  HDNAN4D1 U833 ( .A1(n362), .A2(n363), .A3(n364), .A4(n365), .Z(n356) );
  HDNAN4D1 U832 ( .A1(n358), .A2(n359), .A3(n360), .A4(n361), .Z(n357) );
  HDNAN4D1 U830 ( .A1(n350), .A2(n351), .A3(n352), .A4(n353), .Z(n334) );
  HDNAN4D1 U829 ( .A1(n346), .A2(n347), .A3(n348), .A4(n349), .Z(n335) );
  HDNAN4D1 U828 ( .A1(n342), .A2(n343), .A3(n344), .A4(n345), .Z(n336) );
  HDNAN4D1 U827 ( .A1(n338), .A2(n339), .A3(n340), .A4(n341), .Z(n337) );
  HDAO32DL U40 ( .A1(n201), .A2(n202), .A3(ecl_alu_out_sel_sum_e_l), .B1(n951), 
        .B2(n203), .Z(alu_ecl_zhigh_e) );
  HDADFULD1 addsub_adder_add_24_2_DP_OP_276_5026_1_U2 ( .A(
        byp_alu_rs1_data_e[63]), .B(alu_ecl_adderin2_63_e), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n2), .CO(addsub_cout64_e), .S(
        alu_ecl_adder_out_63_e) );
  HDADFULD1 addsub_adder_add_24_2_DP_OP_276_5026_1_U36 ( .A(
        byp_alu_rs1_data_e[31]), .B(alu_ecl_adderin2_31_e), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n35), .CO(alu_ecl_cout32_e), 
        .S(exu_ifu_brpc_e_31_) );
  HDADFULD1 addsub_adder_add_24_2_DP_OP_276_5026_1_U67 ( .A(
        byp_alu_rs1_data_e[0]), .B(addsub_rs2_data_0), .CI(ecl_alu_cin_e), 
        .CO(addsub_adder_add_24_2_DP_OP_276_5026_1_n65), .S(
        exu_mmu_early_va_e[0]) );
  HDDFFPQ2 invert_d2e_q_reg_0_ ( .D(n940), .CK(rclk), .Q(n7) );
  HDBUFD2 U1109 ( .A(n417), .Z(n939) );
  HDEXNOR2DL U1110 ( .A1(byp_alu_rs2_data_e_l[60]), .A2(addsub_subtract_e[60]), 
        .Z(addsub_rs2_data_60_) );
  HDEXNOR2DL U1111 ( .A1(byp_alu_rs2_data_e_l[5]), .A2(addsub_subtract_e[5]), 
        .Z(addsub_rs2_data_5) );
  HDEXNOR2DL U1112 ( .A1(byp_alu_rs2_data_e_l[13]), .A2(addsub_subtract_e[13]), 
        .Z(addsub_rs2_data_13) );
  HDEXNOR2DL U1113 ( .A1(byp_alu_rs2_data_e_l[26]), .A2(addsub_subtract_e[26]), 
        .Z(addsub_rs2_data_26) );
  HDEXNOR2DL U1114 ( .A1(byp_alu_rs2_data_e_l[35]), .A2(addsub_subtract_e[35]), 
        .Z(addsub_rs2_data_35_) );
  HDEXNOR2DL U1115 ( .A1(byp_alu_rs2_data_e_l[41]), .A2(addsub_subtract_e[41]), 
        .Z(addsub_rs2_data_41_) );
  HDEXNOR2DL U1116 ( .A1(byp_alu_rs2_data_e_l[61]), .A2(addsub_subtract_e[61]), 
        .Z(addsub_rs2_data_61_) );
  HDAOI22D1 U1117 ( .A1(byp_alu_rs1_data_e[43]), .A2(n292), .B1(
        byp_alu_rs1_data_e[42]), .B2(n296), .Z(n930) );
  HDOAI21D1 U1118 ( .A1(byp_alu_rs1_data_e[44]), .A2(addsub_rs2_data_44_), .B(
        n290), .Z(n931) );
  HDOAI21D1 U1119 ( .A1(byp_alu_rs1_data_e[45]), .A2(addsub_rs2_data_45_), .B(
        n293), .Z(n932) );
  HDAOI22D1 U1120 ( .A1(addsub_rs2_data_46_), .A2(n252), .B1(
        byp_alu_rs1_data_e[47]), .B2(n253), .Z(n933) );
  HDNAN4D1 U1121 ( .A1(n930), .A2(n931), .A3(n932), .A4(n933), .Z(n301) );
  HDEXNOR2DL U1122 ( .A1(byp_alu_rs2_data_e_l[6]), .A2(addsub_subtract_e[6]), 
        .Z(addsub_rs2_data_6) );
  HDEXNOR2DL U1123 ( .A1(byp_alu_rs2_data_e_l[27]), .A2(addsub_subtract_e[27]), 
        .Z(addsub_rs2_data_27) );
  HDEXNOR2DL U1124 ( .A1(byp_alu_rs2_data_e_l[36]), .A2(addsub_subtract_e[36]), 
        .Z(addsub_rs2_data_36_) );
  HDEXNOR2DL U1125 ( .A1(byp_alu_rs2_data_e_l[42]), .A2(addsub_subtract_e[42]), 
        .Z(addsub_rs2_data_42_) );
  HDEXNOR2DL U1126 ( .A1(byp_alu_rs2_data_e_l[62]), .A2(addsub_subtract_e[62]), 
        .Z(addsub_rs2_data_62_) );
  HDEXNOR2DL U1127 ( .A1(byp_alu_rs2_data_e_l[0]), .A2(addsub_subtract_e[0]), 
        .Z(addsub_rs2_data_0) );
  HDEXNOR2DL U1128 ( .A1(byp_alu_rs2_data_e_l[7]), .A2(addsub_subtract_e[7]), 
        .Z(addsub_rs2_data_7) );
  HDEXNOR2DL U1129 ( .A1(byp_alu_rs2_data_e_l[28]), .A2(addsub_subtract_e[28]), 
        .Z(addsub_rs2_data_28) );
  HDEXNOR2DL U1130 ( .A1(byp_alu_rs2_data_e_l[37]), .A2(addsub_subtract_e[37]), 
        .Z(addsub_rs2_data_37_) );
  HDEXNOR2DL U1131 ( .A1(byp_alu_rs2_data_e_l[44]), .A2(addsub_subtract_e[44]), 
        .Z(addsub_rs2_data_44_) );
  HDEXNOR2DL U1132 ( .A1(byp_alu_rs2_data_e_l[55]), .A2(addsub_subtract_e[55]), 
        .Z(addsub_rs2_data_55_) );
  HDNOR3DL U1133 ( .A1(byp_alu_rs1_data_e[57]), .A2(addsub_rs2_data_57_), .A3(
        n234), .Z(n934) );
  HDNAN2M1D1 U1134 ( .A1(n144), .A2(n222), .Z(n935) );
  HDOAI31DL U1135 ( .A1(byp_alu_rs1_data_e[61]), .A2(addsub_rs2_data_61_), 
        .A3(n243), .B(n935), .Z(n936) );
  HDOAI33DL U1136 ( .A1(byp_alu_rs1_data_e[59]), .A2(addsub_rs2_data_59_), 
        .A3(n232), .B1(byp_alu_rs1_data_e[58]), .B2(addsub_rs2_data_58_), .B3(
        n233), .Z(n937) );
  HDOAI33DL U1137 ( .A1(byp_alu_rs1_data_e[60]), .A2(addsub_rs2_data_60_), 
        .A3(n242), .B1(byp_alu_rs1_data_e[56]), .B2(addsub_rs2_data_56_), .B3(
        n237), .Z(n938) );
  HDNOR4D1 U1138 ( .A1(n934), .A2(n936), .A3(n937), .A4(n938), .Z(n209) );
  HDEXNOR2DL U1139 ( .A1(byp_alu_rs2_data_e_l[1]), .A2(addsub_subtract_e[1]), 
        .Z(addsub_rs2_data_1) );
  HDEXNOR2DL U1140 ( .A1(byp_alu_rs2_data_e_l[8]), .A2(addsub_subtract_e[8]), 
        .Z(addsub_rs2_data_8) );
  HDEXNOR2DL U1141 ( .A1(byp_alu_rs2_data_e_l[15]), .A2(addsub_subtract_e[15]), 
        .Z(addsub_rs2_data_15) );
  HDEXNOR2DL U1142 ( .A1(byp_alu_rs2_data_e_l[18]), .A2(addsub_subtract_e[18]), 
        .Z(addsub_rs2_data_18) );
  HDEXNOR2DL U1143 ( .A1(byp_alu_rs2_data_e_l[29]), .A2(addsub_subtract_e[29]), 
        .Z(addsub_rs2_data_29) );
  HDEXNOR2DL U1144 ( .A1(byp_alu_rs2_data_e_l[39]), .A2(addsub_subtract_e[39]), 
        .Z(addsub_rs2_data_39_) );
  HDEXNOR2DL U1145 ( .A1(byp_alu_rs2_data_e_l[43]), .A2(addsub_subtract_e[43]), 
        .Z(addsub_rs2_data_43_) );
  HDEXNOR2DL U1146 ( .A1(byp_alu_rs2_data_e_l[46]), .A2(addsub_subtract_e[46]), 
        .Z(addsub_rs2_data_46_) );
  HDEXNOR2DL U1147 ( .A1(byp_alu_rs2_data_e_l[2]), .A2(addsub_subtract_e[2]), 
        .Z(addsub_rs2_data_2) );
  HDEXNOR2DL U1148 ( .A1(byp_alu_rs2_data_e_l[9]), .A2(addsub_subtract_e[9]), 
        .Z(addsub_rs2_data_9) );
  HDEXNOR2DL U1149 ( .A1(byp_alu_rs2_data_e_l[14]), .A2(addsub_subtract_e[14]), 
        .Z(addsub_rs2_data_14) );
  HDEXNOR2DL U1150 ( .A1(byp_alu_rs2_data_e_l[16]), .A2(addsub_subtract_e[16]), 
        .Z(addsub_rs2_data_16) );
  HDEXNOR2DL U1151 ( .A1(byp_alu_rs2_data_e_l[17]), .A2(addsub_subtract_e[17]), 
        .Z(addsub_rs2_data_17) );
  HDEXNOR2DL U1152 ( .A1(byp_alu_rs2_data_e_l[19]), .A2(addsub_subtract_e[19]), 
        .Z(addsub_rs2_data_19) );
  HDEXNOR2DL U1153 ( .A1(byp_alu_rs2_data_e_l[30]), .A2(addsub_subtract_e[30]), 
        .Z(addsub_rs2_data_30) );
  HDEXNOR2DL U1154 ( .A1(byp_alu_rs2_data_e_l[45]), .A2(addsub_subtract_e[45]), 
        .Z(addsub_rs2_data_45_) );
  HDEXNOR2DL U1155 ( .A1(byp_alu_rs2_data_e_l[47]), .A2(addsub_subtract_e[47]), 
        .Z(addsub_rs2_data_47_) );
  HDEXNOR2DL U1156 ( .A1(byp_alu_rs2_data_e_l[31]), .A2(addsub_subtract_e[31]), 
        .Z(alu_ecl_adderin2_31_e) );
  HDEXNOR2DL U1157 ( .A1(byp_alu_rs2_data_e_l[63]), .A2(addsub_subtract_e[63]), 
        .Z(alu_ecl_adderin2_63_e) );
  HDNAN2M1D1 U1158 ( .A1(se), .A2(ifu_exu_invert_d), .Z(n940) );
  HDINVBD4 U1159 ( .A(n7), .Z(invert_e) );
  HDAOI22D1 U1160 ( .A1(n60), .A2(addsub_rs2_data_30), .B1(n63), .B2(
        addsub_rs2_data_29), .Z(n141) );
  HDAOI22D1 U1161 ( .A1(byp_alu_rs1_data_e[15]), .A2(n105), .B1(n104), .B2(
        addsub_rs2_data_16), .Z(n118) );
  HDAOI22D1 U1162 ( .A1(byp_alu_rs1_data_e[58]), .A2(n233), .B1(n232), .B2(
        addsub_rs2_data_59_), .Z(n239) );
  HDAOI22D1 U1163 ( .A1(byp_alu_rs1_data_e[2]), .A2(n50), .B1(n51), .B2(
        addsub_rs2_data_3), .Z(n46) );
  HDAOI22D1 U1164 ( .A1(byp_alu_rs1_data_e[9]), .A2(n41), .B1(n40), .B2(
        addsub_rs2_data_10), .Z(n64) );
  HDOAI21D1 U1165 ( .A1(byp_alu_rs1_data_e[25]), .A2(addsub_rs2_data_25), .B(
        n91), .Z(n132) );
  HDOAI21D1 U1166 ( .A1(byp_alu_rs1_data_e[51]), .A2(addsub_rs2_data_51_), .B(
        n260), .Z(n254) );
  HDOAI33D1 U1167 ( .A1(addsub_rs2_data_1), .A2(byp_alu_rs1_data_e[1]), .A3(
        n52), .B1(addsub_rs2_data_0), .B2(byp_alu_rs1_data_e[0]), .B3(n71), 
        .Z(n79) );
  HDAOI22D1 U1168 ( .A1(byp_alu_rs1_data_e[53]), .A2(n259), .B1(n258), .B2(
        addsub_rs2_data_52_), .Z(n255) );
  HDAOI22D1 U1169 ( .A1(n236), .A2(addsub_rs2_data_55_), .B1(n235), .B2(
        addsub_rs2_data_54_), .Z(n256) );
  HDAOI22D1 U1170 ( .A1(byp_alu_rs1_data_e[52]), .A2(n258), .B1(n259), .B2(
        addsub_rs2_data_53_), .Z(n257) );
  HDAOI22D1 U1171 ( .A1(byp_alu_rs1_data_e[21]), .A2(n95), .B1(n94), .B2(
        addsub_rs2_data_22), .Z(n131) );
  HDAOI22D1 U1172 ( .A1(n250), .A2(addsub_rs2_data_49_), .B1(n249), .B2(
        addsub_rs2_data_48_), .Z(n245) );
  HDAOI22D1 U1173 ( .A1(byp_alu_rs1_data_e[46]), .A2(n252), .B1(n253), .B2(
        addsub_rs2_data_47_), .Z(n246) );
  HDOAI21D1 U1174 ( .A1(byp_alu_rs1_data_e[50]), .A2(addsub_rs2_data_50_), .B(
        n251), .Z(n247) );
  HDAOI22D1 U1175 ( .A1(n92), .A2(addsub_rs2_data_24), .B1(n96), .B2(
        addsub_rs2_data_23), .Z(n130) );
  HDOAI21D1 U1176 ( .A1(byp_alu_rs1_data_e[26]), .A2(addsub_rs2_data_26), .B(
        n93), .Z(n139) );
  HDAOI22D1 U1177 ( .A1(byp_alu_rs1_data_e[28]), .A2(n61), .B1(n62), .B2(
        addsub_rs2_data_27), .Z(n140) );
  HDOAI33D1 U1178 ( .A1(addsub_rs2_data_19), .A2(byp_alu_rs1_data_e[19]), .A3(
        n97), .B1(addsub_rs2_data_18), .B2(byp_alu_rs1_data_e[18]), .B3(n98), 
        .Z(n87) );
  HDAOI22D1 U1179 ( .A1(byp_alu_rs1_data_e[59]), .A2(n232), .B1(n233), .B2(
        addsub_rs2_data_58_), .Z(n231) );
  HDOAI21D1 U1180 ( .A1(byp_alu_rs1_data_e[57]), .A2(addsub_rs2_data_57_), .B(
        n234), .Z(n230) );
  HDAOI22D1 U1181 ( .A1(byp_alu_rs1_data_e[27]), .A2(n62), .B1(n61), .B2(
        addsub_rs2_data_28), .Z(n142) );
  HDOAI21D1 U1182 ( .A1(byp_alu_rs1_data_e[56]), .A2(addsub_rs2_data_56_), .B(
        n237), .Z(n228) );
  HDAOI22D1 U1183 ( .A1(n243), .A2(addsub_rs2_data_61_), .B1(n242), .B2(
        addsub_rs2_data_60_), .Z(n238) );
  HDOAI33D1 U1184 ( .A1(addsub_rs2_data_13), .A2(byp_alu_rs1_data_e[13]), .A3(
        n69), .B1(addsub_rs2_data_12), .B2(byp_alu_rs1_data_e[12]), .B3(n68), 
        .Z(n100) );
  HDOAI21D1 U1185 ( .A1(byp_alu_rs1_data_e[62]), .A2(addsub_rs2_data_62_), .B(
        n244), .Z(n240) );
  HDOAI33D1 U1186 ( .A1(addsub_rs2_data_15), .A2(byp_alu_rs1_data_e[15]), .A3(
        n105), .B1(addsub_rs2_data_17), .B2(byp_alu_rs1_data_e[17]), .B3(n106), 
        .Z(n101) );
  HDAOI22D1 U1187 ( .A1(n220), .A2(addsub_rs2_data_36_), .B1(n216), .B2(
        addsub_rs2_data_37_), .Z(n326) );
  HDOAI21D1 U1188 ( .A1(byp_alu_rs1_data_e[14]), .A2(addsub_rs2_data_14), .B(
        n109), .Z(n115) );
  HDAOI22D1 U1189 ( .A1(byp_alu_rs1_data_e[22]), .A2(n94), .B1(n95), .B2(
        addsub_rs2_data_21), .Z(n125) );
  HDAOI22D1 U1190 ( .A1(n296), .A2(addsub_rs2_data_42_), .B1(n292), .B2(
        addsub_rs2_data_43_), .Z(n319) );
  HDAOI22D1 U1191 ( .A1(byp_alu_rs1_data_e[37]), .A2(n216), .B1(n297), .B2(
        addsub_rs2_data_38_), .Z(n328) );
  HDOAI21D1 U1192 ( .A1(byp_alu_rs1_data_e[7]), .A2(addsub_rs2_data_7), .B(n42), .Z(n36) );
  HDAOI22D1 U1193 ( .A1(byp_alu_rs1_data_e[34]), .A2(n219), .B1(n218), .B2(
        addsub_rs2_data_35_), .Z(n325) );
  HDAOI22D1 U1194 ( .A1(byp_alu_rs1_data_e[5]), .A2(n43), .B1(n44), .B2(
        addsub_rs2_data_6), .Z(n35) );
  HDAOI22D1 U1195 ( .A1(byp_alu_rs1_data_e[40]), .A2(n295), .B1(n294), .B2(
        addsub_rs2_data_41_), .Z(n318) );
  HDAOI22D1 U1196 ( .A1(n39), .A2(addsub_rs2_data_8), .B1(n41), .B2(
        addsub_rs2_data_9), .Z(n37) );
  HDAOI22D1 U1197 ( .A1(n223), .A2(addsub_rs2_data_33_), .B1(n219), .B2(
        addsub_rs2_data_34_), .Z(n299) );
  HDAOI22D1 U1198 ( .A1(byp_alu_rs1_data_e[31]), .A2(n222), .B1(n221), .B2(
        addsub_rs2_data_32_), .Z(n298) );
  HDAOI22D1 U1199 ( .A1(n217), .A2(addsub_rs2_data_39_), .B1(n295), .B2(
        addsub_rs2_data_40_), .Z(n316) );
  HDOAI21D1 U1200 ( .A1(byp_alu_rs1_data_e[20]), .A2(addsub_rs2_data_20), .B(
        n103), .Z(n124) );
  HDAOI22D1 U1201 ( .A1(n43), .A2(addsub_rs2_data_5), .B1(n49), .B2(
        addsub_rs2_data_4), .Z(n47) );
  HDBUFD2 U1202 ( .A(n450), .Z(n941) );
  HDADFULDL U1203 ( .A(byp_alu_rs1_data_e[2]), .B(addsub_rs2_data_2), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n64), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n63), .S(exu_mmu_early_va_e[2])
         );
  HDOR3DL U1204 ( .A1(byp_alu_rs1_data_e[2]), .A2(n50), .A3(addsub_rs2_data_2), 
        .Z(n84) );
  HDADFULDL U1205 ( .A(byp_alu_rs1_data_e[55]), .B(addsub_rs2_data_55_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n10), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n9), .S(adder_out[55]) );
  HDOR3DL U1206 ( .A1(byp_alu_rs1_data_e[55]), .A2(n236), .A3(
        addsub_rs2_data_55_), .Z(n274) );
  HDADFULDL U1207 ( .A(byp_alu_rs1_data_e[57]), .B(addsub_rs2_data_57_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n8), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n7), .S(adder_out[57]) );
  HDADFULDL U1208 ( .A(byp_alu_rs1_data_e[1]), .B(addsub_rs2_data_1), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n65), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n64), .S(exu_mmu_early_va_e[1])
         );
  HDAOI222DL U1209 ( .A1(n71), .A2(n72), .B1(n50), .B2(addsub_rs2_data_2), 
        .C1(n52), .C2(addsub_rs2_data_1), .Z(n55) );
  HDADFULDL U1210 ( .A(byp_alu_rs1_data_e[61]), .B(addsub_rs2_data_61_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n4), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n3), .S(adder_out[61]) );
  HDADFULDL U1211 ( .A(byp_alu_rs1_data_e[47]), .B(addsub_rs2_data_47_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n18), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n17), .S(exu_ifu_brpc_e[47]) );
  HDADFULDL U1212 ( .A(byp_alu_rs1_data_e[43]), .B(addsub_rs2_data_43_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n22), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n21), .S(exu_ifu_brpc_e[43]) );
  HDADFULDL U1213 ( .A(byp_alu_rs1_data_e[41]), .B(addsub_rs2_data_41_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n24), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n23), .S(exu_ifu_brpc_e[41]) );
  HDADFULDL U1214 ( .A(byp_alu_rs1_data_e[37]), .B(addsub_rs2_data_37_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n28), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n27), .S(exu_ifu_brpc_e[37]) );
  HDADFULDL U1215 ( .A(byp_alu_rs1_data_e[35]), .B(addsub_rs2_data_35_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n30), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n29), .S(exu_ifu_brpc_e[35]) );
  HDADFULDL U1216 ( .A(byp_alu_rs1_data_e[27]), .B(addsub_rs2_data_27), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n39), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n38), .S(exu_ifu_brpc_e[27]) );
  HDADFULDL U1217 ( .A(byp_alu_rs1_data_e[21]), .B(addsub_rs2_data_21), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n45), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n44), .S(exu_ifu_brpc_e[21]) );
  HDADFULDL U1218 ( .A(byp_alu_rs1_data_e[15]), .B(addsub_rs2_data_15), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n51), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n50), .S(exu_ifu_brpc_e[15]) );
  HDAOI22DL U1219 ( .A1(byp_alu_rs1_data_e[16]), .A2(n104), .B1(n105), .B2(
        addsub_rs2_data_15), .Z(n116) );
  HDADFULDL U1220 ( .A(byp_alu_rs1_data_e[13]), .B(addsub_rs2_data_13), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n53), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n52), .S(exu_ifu_brpc_e[13]) );
  HDAOI22DL U1221 ( .A1(byp_alu_rs1_data_e[12]), .A2(n68), .B1(n69), .B2(
        addsub_rs2_data_13), .Z(n67) );
  HDADFULDL U1222 ( .A(byp_alu_rs1_data_e[9]), .B(addsub_rs2_data_9), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n57), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n56), .S(exu_lsu_early_va_e[9])
         );
  HDADFULDL U1223 ( .A(byp_alu_rs1_data_e[3]), .B(addsub_rs2_data_3), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n63), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n62), .S(exu_lsu_early_va_e[3])
         );
  HDADFULDL U1224 ( .A(byp_alu_rs1_data_e[60]), .B(addsub_rs2_data_60_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n5), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n4), .S(adder_out[60]) );
  HDADFULDL U1225 ( .A(byp_alu_rs1_data_e[59]), .B(addsub_rs2_data_59_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n6), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n5), .S(adder_out[59]) );
  HDADFULDL U1226 ( .A(byp_alu_rs1_data_e[54]), .B(addsub_rs2_data_54_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n11), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n10), .S(adder_out[54]) );
  HDADFULDL U1227 ( .A(byp_alu_rs1_data_e[53]), .B(addsub_rs2_data_53_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n12), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n11), .S(adder_out[53]) );
  HDADFULDL U1228 ( .A(byp_alu_rs1_data_e[48]), .B(addsub_rs2_data_48_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n17), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n16), .S(adder_out[48]) );
  HDADFULDL U1229 ( .A(byp_alu_rs1_data_e[42]), .B(addsub_rs2_data_42_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n23), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n22), .S(exu_ifu_brpc_e[42]) );
  HDADFULDL U1230 ( .A(byp_alu_rs1_data_e[36]), .B(addsub_rs2_data_36_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n29), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n28), .S(exu_ifu_brpc_e[36]) );
  HDADFULDL U1231 ( .A(byp_alu_rs1_data_e[30]), .B(addsub_rs2_data_30), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n36), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n35), .S(exu_ifu_brpc_e[30]) );
  HDADFULDL U1232 ( .A(byp_alu_rs1_data_e[8]), .B(addsub_rs2_data_8), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n58), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n57), .S(exu_lsu_early_va_e[8])
         );
  HDADFULDL U1233 ( .A(byp_alu_rs1_data_e[49]), .B(addsub_rs2_data_49_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n16), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n15), .S(adder_out[49]) );
  HDADFULDL U1234 ( .A(byp_alu_rs1_data_e[45]), .B(addsub_rs2_data_45_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n20), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n19), .S(exu_ifu_brpc_e[45]) );
  HDOAI33DL U1235 ( .A1(addsub_rs2_data_43_), .A2(byp_alu_rs1_data_e[43]), 
        .A3(n292), .B1(addsub_rs2_data_45_), .B2(byp_alu_rs1_data_e[45]), .B3(
        n293), .Z(n288) );
  HDADFULDL U1236 ( .A(byp_alu_rs1_data_e[44]), .B(addsub_rs2_data_44_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n21), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n20), .S(exu_ifu_brpc_e[44]) );
  HDOAI33DL U1237 ( .A1(addsub_rs2_data_48_), .A2(byp_alu_rs1_data_e[48]), 
        .A3(n249), .B1(addsub_rs2_data_44_), .B2(byp_alu_rs1_data_e[44]), .B3(
        n290), .Z(n289) );
  HDADFULDL U1238 ( .A(byp_alu_rs1_data_e[40]), .B(addsub_rs2_data_40_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n25), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n24), .S(exu_ifu_brpc_e[40]) );
  HDOAI33DL U1239 ( .A1(addsub_rs2_data_41_), .A2(byp_alu_rs1_data_e[41]), 
        .A3(n294), .B1(addsub_rs2_data_40_), .B2(byp_alu_rs1_data_e[40]), .B3(
        n295), .Z(n287) );
  HDADFULDL U1240 ( .A(byp_alu_rs1_data_e[38]), .B(addsub_rs2_data_38_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n27), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n26), .S(exu_ifu_brpc_e[38]) );
  HDOAI33DL U1241 ( .A1(addsub_rs2_data_42_), .A2(byp_alu_rs1_data_e[42]), 
        .A3(n296), .B1(addsub_rs2_data_38_), .B2(byp_alu_rs1_data_e[38]), .B3(
        n297), .Z(n286) );
  HDADFULDL U1242 ( .A(byp_alu_rs1_data_e[34]), .B(addsub_rs2_data_34_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n31), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n30), .S(exu_ifu_brpc_e[34]) );
  HDOAI33DL U1243 ( .A1(addsub_rs2_data_35_), .A2(byp_alu_rs1_data_e[35]), 
        .A3(n218), .B1(addsub_rs2_data_34_), .B2(byp_alu_rs1_data_e[34]), .B3(
        n219), .Z(n214) );
  HDADFULDL U1244 ( .A(byp_alu_rs1_data_e[32]), .B(addsub_rs2_data_32_), .CI(
        alu_ecl_cout32_e), .CO(addsub_adder_add_24_2_DP_OP_276_5026_1_n32), 
        .S(exu_ifu_brpc_e[32]) );
  HDOAI33DL U1245 ( .A1(addsub_rs2_data_36_), .A2(byp_alu_rs1_data_e[36]), 
        .A3(n220), .B1(addsub_rs2_data_32_), .B2(byp_alu_rs1_data_e[32]), .B3(
        n221), .Z(n213) );
  HDADFULDL U1246 ( .A(byp_alu_rs1_data_e[29]), .B(addsub_rs2_data_29), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n37), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n36), .S(exu_ifu_brpc_e[29]) );
  HDOAI33DL U1247 ( .A1(addsub_rs2_data_27), .A2(byp_alu_rs1_data_e[27]), .A3(
        n62), .B1(addsub_rs2_data_29), .B2(byp_alu_rs1_data_e[29]), .B3(n63), 
        .Z(n58) );
  HDADFULDL U1248 ( .A(byp_alu_rs1_data_e[28]), .B(addsub_rs2_data_28), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n38), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n37), .S(exu_ifu_brpc_e[28]) );
  HDOAI33DL U1249 ( .A1(addsub_rs2_data_30), .A2(byp_alu_rs1_data_e[30]), .A3(
        n60), .B1(addsub_rs2_data_28), .B2(byp_alu_rs1_data_e[28]), .B3(n61), 
        .Z(n59) );
  HDADFULDL U1250 ( .A(byp_alu_rs1_data_e[23]), .B(addsub_rs2_data_23), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n43), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n42), .S(exu_ifu_brpc_e[23]) );
  HDOAI33DL U1251 ( .A1(addsub_rs2_data_21), .A2(byp_alu_rs1_data_e[21]), .A3(
        n95), .B1(addsub_rs2_data_23), .B2(byp_alu_rs1_data_e[23]), .B3(n96), 
        .Z(n88) );
  HDADFULDL U1252 ( .A(byp_alu_rs1_data_e[22]), .B(addsub_rs2_data_22), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n44), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n43), .S(exu_ifu_brpc_e[22]) );
  HDADFULDL U1253 ( .A(byp_alu_rs1_data_e[17]), .B(addsub_rs2_data_17), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n49), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n48), .S(exu_ifu_brpc_e[17]) );
  HDADFULDL U1254 ( .A(byp_alu_rs1_data_e[16]), .B(addsub_rs2_data_16), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n50), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n49), .S(exu_ifu_brpc_e[16]) );
  HDADFULDL U1255 ( .A(byp_alu_rs1_data_e[12]), .B(addsub_rs2_data_12), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n54), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n53), .S(exu_ifu_brpc_e[12]) );
  HDADFULDL U1256 ( .A(byp_alu_rs1_data_e[10]), .B(addsub_rs2_data_10), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n56), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n55), .S(exu_lsu_early_va_e[10]) );
  HDADFULDL U1257 ( .A(byp_alu_rs1_data_e[6]), .B(addsub_rs2_data_6), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n60), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n59), .S(exu_lsu_early_va_e[6])
         );
  HDADFULDL U1258 ( .A(byp_alu_rs1_data_e[4]), .B(addsub_rs2_data_4), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n62), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n61), .S(exu_lsu_early_va_e[4])
         );
  HDOAI33DL U1259 ( .A1(addsub_rs2_data_8), .A2(byp_alu_rs1_data_e[8]), .A3(
        n39), .B1(addsub_rs2_data_4), .B2(byp_alu_rs1_data_e[4]), .B3(n49), 
        .Z(n150) );
  HDADFULDL U1260 ( .A(byp_alu_rs1_data_e[58]), .B(addsub_rs2_data_58_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n7), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n6), .S(adder_out[58]) );
  HDADFULDL U1261 ( .A(byp_alu_rs1_data_e[52]), .B(addsub_rs2_data_52_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n13), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n12), .S(adder_out[52]) );
  HDOAI33DL U1262 ( .A1(addsub_rs2_data_53_), .A2(byp_alu_rs1_data_e[53]), 
        .A3(n259), .B1(addsub_rs2_data_52_), .B2(byp_alu_rs1_data_e[52]), .B3(
        n258), .Z(n279) );
  HDADFULDL U1263 ( .A(byp_alu_rs1_data_e[46]), .B(addsub_rs2_data_46_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n19), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n18), .S(exu_ifu_brpc_e[46]) );
  HDOAI33DL U1264 ( .A1(addsub_rs2_data_47_), .A2(byp_alu_rs1_data_e[47]), 
        .A3(n253), .B1(addsub_rs2_data_46_), .B2(byp_alu_rs1_data_e[46]), .B3(
        n252), .Z(n276) );
  HDADFULDL U1265 ( .A(byp_alu_rs1_data_e[39]), .B(addsub_rs2_data_39_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n26), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n25), .S(exu_ifu_brpc_e[39]) );
  HDOAI33DL U1266 ( .A1(addsub_rs2_data_37_), .A2(byp_alu_rs1_data_e[37]), 
        .A3(n216), .B1(addsub_rs2_data_39_), .B2(byp_alu_rs1_data_e[39]), .B3(
        n217), .Z(n215) );
  HDADFULDL U1267 ( .A(byp_alu_rs1_data_e[33]), .B(addsub_rs2_data_33_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n32), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n31), .S(exu_ifu_brpc_e[33]) );
  HDOAI33DL U1268 ( .A1(alu_ecl_adderin2_31_e), .A2(byp_alu_rs1_data_e[31]), 
        .A3(n222), .B1(addsub_rs2_data_33_), .B2(byp_alu_rs1_data_e[33]), .B3(
        n223), .Z(n212) );
  HDADFULDL U1269 ( .A(byp_alu_rs1_data_e[24]), .B(addsub_rs2_data_24), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n42), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n41), .S(exu_ifu_brpc_e[24]) );
  HDADFULDL U1270 ( .A(byp_alu_rs1_data_e[18]), .B(addsub_rs2_data_18), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n48), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n47), .S(exu_ifu_brpc_e[18]) );
  HDAOI22DL U1271 ( .A1(n98), .A2(addsub_rs2_data_18), .B1(n106), .B2(
        addsub_rs2_data_17), .Z(n117) );
  HDADFULDL U1272 ( .A(byp_alu_rs1_data_e[11]), .B(addsub_rs2_data_11), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n55), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n54), .S(exu_ifu_brpc_e[11]) );
  HDAOI22DL U1273 ( .A1(n70), .A2(addsub_rs2_data_11), .B1(n68), .B2(
        addsub_rs2_data_12), .Z(n65) );
  HDOAI33DL U1274 ( .A1(addsub_rs2_data_9), .A2(byp_alu_rs1_data_e[9]), .A3(
        n41), .B1(addsub_rs2_data_11), .B2(byp_alu_rs1_data_e[11]), .B3(n70), 
        .Z(n152) );
  HDADFULDL U1275 ( .A(byp_alu_rs1_data_e[5]), .B(addsub_rs2_data_5), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n61), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n60), .S(exu_lsu_early_va_e[5])
         );
  HDOAI33DL U1276 ( .A1(addsub_rs2_data_3), .A2(byp_alu_rs1_data_e[3]), .A3(
        n51), .B1(addsub_rs2_data_5), .B2(byp_alu_rs1_data_e[5]), .B3(n43), 
        .Z(n149) );
  HDADFULDL U1277 ( .A(byp_alu_rs1_data_e[26]), .B(addsub_rs2_data_26), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n40), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n39), .S(exu_ifu_brpc_e[26]) );
  HDOAI33DL U1278 ( .A1(addsub_rs2_data_26), .A2(byp_alu_rs1_data_e[26]), .A3(
        n93), .B1(addsub_rs2_data_22), .B2(byp_alu_rs1_data_e[22]), .B3(n94), 
        .Z(n89) );
  HDADFULDL U1279 ( .A(byp_alu_rs1_data_e[25]), .B(addsub_rs2_data_25), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n41), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n40), .S(exu_ifu_brpc_e[25]) );
  HDOAI33DL U1280 ( .A1(addsub_rs2_data_25), .A2(byp_alu_rs1_data_e[25]), .A3(
        n91), .B1(addsub_rs2_data_24), .B2(byp_alu_rs1_data_e[24]), .B3(n92), 
        .Z(n90) );
  HDADFULDL U1281 ( .A(byp_alu_rs1_data_e[20]), .B(addsub_rs2_data_20), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n46), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n45), .S(exu_ifu_brpc_e[20]) );
  HDOAI33DL U1282 ( .A1(addsub_rs2_data_20), .A2(byp_alu_rs1_data_e[20]), .A3(
        n103), .B1(addsub_rs2_data_16), .B2(byp_alu_rs1_data_e[16]), .B3(n104), 
        .Z(n102) );
  HDADFULDL U1283 ( .A(byp_alu_rs1_data_e[19]), .B(addsub_rs2_data_19), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n47), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n46), .S(exu_ifu_brpc_e[19]) );
  HDOAI21DL U1284 ( .A1(byp_alu_rs1_data_e[19]), .A2(addsub_rs2_data_19), .B(
        n97), .Z(n122) );
  HDADFULDL U1285 ( .A(byp_alu_rs1_data_e[14]), .B(addsub_rs2_data_14), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n52), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n51), .S(exu_ifu_brpc_e[14]) );
  HDOAI33DL U1286 ( .A1(addsub_rs2_data_14), .A2(byp_alu_rs1_data_e[14]), .A3(
        n109), .B1(addsub_rs2_data_10), .B2(byp_alu_rs1_data_e[10]), .B3(n40), 
        .Z(n99) );
  HDADFULDL U1287 ( .A(byp_alu_rs1_data_e[7]), .B(addsub_rs2_data_7), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n59), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n58), .S(exu_lsu_early_va_e[7])
         );
  HDOAI33DL U1288 ( .A1(addsub_rs2_data_7), .A2(byp_alu_rs1_data_e[7]), .A3(
        n42), .B1(addsub_rs2_data_6), .B2(byp_alu_rs1_data_e[6]), .B3(n44), 
        .Z(n151) );
  HDADFULDL U1289 ( .A(byp_alu_rs1_data_e[56]), .B(addsub_rs2_data_56_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n9), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n8), .S(adder_out[56]) );
  HDADFULDL U1290 ( .A(byp_alu_rs1_data_e[51]), .B(addsub_rs2_data_51_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n14), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n13), .S(adder_out[51]) );
  HDOAI33DL U1291 ( .A1(addsub_rs2_data_49_), .A2(byp_alu_rs1_data_e[49]), 
        .A3(n250), .B1(addsub_rs2_data_51_), .B2(byp_alu_rs1_data_e[51]), .B3(
        n260), .Z(n277) );
  HDADFULDL U1292 ( .A(byp_alu_rs1_data_e[50]), .B(addsub_rs2_data_50_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n15), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n14), .S(adder_out[50]) );
  HDOAI33DL U1293 ( .A1(addsub_rs2_data_54_), .A2(byp_alu_rs1_data_e[54]), 
        .A3(n235), .B1(addsub_rs2_data_50_), .B2(byp_alu_rs1_data_e[50]), .B3(
        n251), .Z(n278) );
  HDADFULDL U1294 ( .A(byp_alu_rs1_data_e[62]), .B(addsub_rs2_data_62_), .CI(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n3), .CO(
        addsub_adder_add_24_2_DP_OP_276_5026_1_n2), .S(adder_out[62]) );
  HDOAI31DL U1295 ( .A1(addsub_rs2_data_62_), .A2(byp_alu_rs1_data_e[62]), 
        .A3(n244), .B(n303), .Z(n302) );
  HDNOR2DL U1296 ( .A1(byp_alu_rs2_data_e_l[47]), .A2(n941), .Z(n577) );
  HDNOR2DL U1297 ( .A1(byp_alu_rs2_data_e_l[54]), .A2(n941), .Z(n521) );
  HDNOR2DL U1298 ( .A1(byp_alu_rs2_data_e_l[41]), .A2(n941), .Z(n619) );
  HDNOR2DL U1299 ( .A1(byp_alu_rs2_data_e_l[40]), .A2(n941), .Z(n626) );
  HDNOR2DL U1300 ( .A1(byp_alu_rs2_data_e_l[39]), .A2(n941), .Z(n640) );
  HDNOR2DL U1301 ( .A1(byp_alu_rs2_data_e_l[46]), .A2(n941), .Z(n584) );
  HDNOR2DL U1302 ( .A1(byp_alu_rs2_data_e_l[45]), .A2(n941), .Z(n591) );
  HDNOR2DL U1303 ( .A1(byp_alu_rs2_data_e_l[44]), .A2(n941), .Z(n598) );
  HDNOR2DL U1304 ( .A1(byp_alu_rs2_data_e_l[43]), .A2(n941), .Z(n605) );
  HDNOR2DL U1305 ( .A1(byp_alu_rs2_data_e_l[34]), .A2(n941), .Z(n675) );
  HDNOR2DL U1306 ( .A1(byp_alu_rs2_data_e_l[32]), .A2(n941), .Z(n689) );
  HDNOR2DL U1307 ( .A1(byp_alu_rs2_data_e_l[38]), .A2(n941), .Z(n647) );
  HDNOR2DL U1308 ( .A1(byp_alu_rs2_data_e_l[37]), .A2(n941), .Z(n654) );
  HDNOR2DL U1309 ( .A1(byp_alu_rs2_data_e_l[36]), .A2(n941), .Z(n661) );
  HDNOR2DL U1310 ( .A1(byp_alu_rs2_data_e_l[35]), .A2(n941), .Z(n668) );
  HDNOR2DL U1311 ( .A1(byp_alu_rs2_data_e_l[58]), .A2(n941), .Z(n493) );
  HDNOR2DL U1312 ( .A1(byp_alu_rs2_data_e_l[57]), .A2(n941), .Z(n500) );
  HDNOR2DL U1313 ( .A1(byp_alu_rs2_data_e_l[56]), .A2(n941), .Z(n507) );
  HDNOR2DL U1314 ( .A1(byp_alu_rs2_data_e_l[53]), .A2(n941), .Z(n528) );
  HDNOR2DL U1315 ( .A1(byp_alu_rs2_data_e_l[42]), .A2(n941), .Z(n612) );
  HDNOR2DL U1316 ( .A1(byp_alu_rs2_data_e_l[55]), .A2(n941), .Z(n514) );
  HDNOR2DL U1317 ( .A1(byp_alu_rs2_data_e_l[50]), .A2(n941), .Z(n549) );
  HDNOR2DL U1318 ( .A1(byp_alu_rs2_data_e_l[49]), .A2(n941), .Z(n563) );
  HDINVBD2 U1319 ( .A(ecl_alu_log_sel_move_e), .Z(n422) );
  HDINVBD2 U1320 ( .A(ecl_alu_out_sel_rs3_e_l), .Z(n417) );
  HDINVD8 U1321 ( .A(n940), .Z(n953) );
  HDINVD1 U1322 ( .A(ecl_alu_out_sel_shift_e_l), .Z(n942) );
  HDINVD1 U1323 ( .A(ecl_alu_out_sel_sum_e_l), .Z(n948) );
  HDINVD1 U1324 ( .A(ecl_alu_out_sel_shift_e_l), .Z(n943) );
  HDINVD1 U1325 ( .A(ecl_alu_out_sel_sum_e_l), .Z(n949) );
  HDINVD1 U1326 ( .A(ecl_alu_out_sel_shift_e_l), .Z(n944) );
  HDINVD1 U1327 ( .A(ecl_alu_out_sel_sum_e_l), .Z(n950) );
  HDINVD1 U1328 ( .A(ecl_alu_out_sel_shift_e_l), .Z(n945) );
  HDINVD1 U1329 ( .A(ecl_alu_out_sel_sum_e_l), .Z(n951) );
  HDINVD1 U1330 ( .A(ecl_alu_out_sel_sum_e_l), .Z(n952) );
  HDINVD1 U1331 ( .A(ecl_alu_out_sel_shift_e_l), .Z(n946) );
  HDINVD2 U1332 ( .A(ecl_alu_out_sel_sum_e_l), .Z(n30) );
  HDINVD1 U1333 ( .A(ecl_alu_out_sel_shift_e_l), .Z(n947) );
  HDINVD2 U1334 ( .A(invert_e), .Z(n956) );
  HDINVD2 U1335 ( .A(invert_e), .Z(n955) );
  HDINVD1 U1336 ( .A(ecl_alu_log_sel_or_e), .Z(n966) );
  HDINVD1 U1337 ( .A(ecl_alu_log_sel_xor_e), .Z(n959) );
  HDINVD1 U1338 ( .A(ecl_alu_log_sel_xor_e), .Z(n962) );
  HDINVD1 U1339 ( .A(ecl_alu_log_sel_or_e), .Z(n968) );
  HDINVD1 U1340 ( .A(ecl_alu_log_sel_xor_e), .Z(n961) );
  HDINVD1 U1341 ( .A(ecl_alu_log_sel_or_e), .Z(n967) );
  HDINVD1 U1342 ( .A(ecl_alu_log_sel_xor_e), .Z(n960) );
  HDINVD1 U1343 ( .A(ecl_alu_log_sel_or_e), .Z(n965) );
  HDINVD1 U1344 ( .A(ecl_alu_log_sel_xor_e), .Z(n958) );
  HDINVD1 U1345 ( .A(ecl_alu_log_sel_or_e), .Z(n964) );
  HDINVD1 U1346 ( .A(ecl_alu_log_sel_xor_e), .Z(n957) );
  HDINVD1 U1347 ( .A(ecl_alu_log_sel_or_e), .Z(n963) );
  HDINVD1 U1348 ( .A(n7), .Z(n954) );
endmodule

