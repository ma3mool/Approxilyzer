
module sparc_exu ( alu_byp_rd_data_e, byp_alu_rs1_data_e, byp_alu_rs2_data_e, 
        ecl_alu_cin_e, ifu_exu_invert_d, ecl_alu_log_sel_and_e, 
        ecl_alu_log_sel_or_e, ecl_alu_log_sel_xor_e, ecl_alu_log_sel_move_e, 
        ecl_alu_out_sel_sum_e_l, ecl_alu_out_sel_shift_e_l, 
        ecl_alu_out_sel_logic_e_l, ecl_alu_sethi_inst_e, ecl_shft_op32_e, 
        ecl_shft_shift4_e, ecl_shft_shift1_e, ecl_shft_enshift_e_l, 
        ecl_shft_extendbit_e, ecl_shft_extend32bit_e_l, ecl_shft_lshift_e_l );
  output [63:0] alu_byp_rd_data_e;
  input [63:0] byp_alu_rs1_data_e;
  input [63:0] byp_alu_rs2_data_e;
  input [3:0] ecl_shft_shift4_e;
  input [3:0] ecl_shft_shift1_e;
  input ecl_alu_cin_e, ifu_exu_invert_d, ecl_alu_log_sel_and_e,
         ecl_alu_log_sel_or_e, ecl_alu_log_sel_xor_e, ecl_alu_log_sel_move_e,
         ecl_alu_out_sel_sum_e_l, ecl_alu_out_sel_shift_e_l,
         ecl_alu_out_sel_logic_e_l, ecl_alu_sethi_inst_e, ecl_shft_op32_e,
         ecl_shft_enshift_e_l, ecl_shft_extendbit_e, ecl_shft_extend32bit_e_l,
         ecl_shft_lshift_e_l;
  wire   alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I2_30_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I2_29_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I2_24_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I2_22_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I2_21_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I2_20_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_29_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_28_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_27_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_26_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_25_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_24_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_23_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_22_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_21_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_19_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_18_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_17_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_15_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_14_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_13_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_12_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_11_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_8_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_7_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_5_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_4_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_3_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n1010,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n1009,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n1006,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n1003,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n1002,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n1000,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n999,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n998,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n997,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n996,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n995,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n992,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n990,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n989,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n985,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n984,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n983,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n982,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n981,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n980,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n977,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n976,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n966,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n961,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n959,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n954,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n953,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n951,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n944,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n938,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n936,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n935,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n933,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n926,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n917,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n916,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n915,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n906,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n905,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n904,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n903,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n902,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n896,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n895,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n894,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n893,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n892,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n886,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n885,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n882,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n881,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n880,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n873,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n872,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n871,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n870,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n869,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n866,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n863,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n862,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n861,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n860,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n855,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n854,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n852,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n851,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n850,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n849,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n848,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n847,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n845,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n843,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n839,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n837,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n828,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n826,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n816,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n813,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n804,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n803,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n802,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n801,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n800,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n799,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n798,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n796,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n793,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n792,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n787,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n777,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n776,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n775,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n774,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n773,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n772,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n766,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n764,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n761,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n752,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n751,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n747,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n746,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n744,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n742,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n739,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n738,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n735,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n726,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n725,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n724,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n723,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n722,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n721,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n720,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n715,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n714,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n713,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n712,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n711,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n710,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n709,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n708,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n707,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n700,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n699,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n698,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n697,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n696,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n695,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n694,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n692,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n689,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n688,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n687,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n686,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n685,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n684,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n683,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n682,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n681,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n676,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n674,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n673,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n672,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n671,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n670,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n669,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n668,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n665,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n663,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n662,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n661,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n660,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n659,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n658,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n657,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n652,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n651,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n649,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n647,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n646,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n645,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n644,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n643,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n642,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n640,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n638,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n636,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n632,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n624,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n620,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n619,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n618,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n617,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n616,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n615,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n614,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n613,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n611,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n609,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n608,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n607,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n606,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n604,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n603,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n602,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n601,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n600,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n599,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n598,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n597,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n596,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n595,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n593,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n591,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n589,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n587,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n583,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n579,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n577,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n575,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n571,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n569,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n565,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n561,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n560,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n544,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n532,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n531,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n515,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n514,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n510,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n508,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n506,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n505,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n499,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n498,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n491,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n481,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n480,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n476,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n474,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n472,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n471,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n465,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n464,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n447,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n446,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n442,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n437,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n435,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n432,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n431,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n430,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n429,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n426,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n423,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n412,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n408,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n404,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n403,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n397,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n396,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n395,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n379,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n370,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n369,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n366,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n364,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n363,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n362,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n361,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n355,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n345,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n344,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n340,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n338,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n332,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n331,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n330,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n329,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n328,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n327,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n321,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n311,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n310,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n306,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n304,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n302,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n301,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n299,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n298,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n297,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n290,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n287,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n277,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n276,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n272,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n270,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n268,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n267,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n262,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n261,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n260,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n259,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n258,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n257,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n256,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n253,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n243,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n242,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n238,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n236,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n234,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n233,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n228,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n227,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n226,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n225,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n219,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n209,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n208,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n204,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n202,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n196,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n195,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n193,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n192,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n191,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n185,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n175,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n174,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n170,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n168,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n166,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n165,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n164,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n163,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n162,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n161,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n159,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n158,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n157,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n141,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n140,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n136,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n128,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n127,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n126,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n125,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n123,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n121,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n120,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n117,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n107,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n106,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n102,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n97,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n96,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n95,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n94,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n93,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n91,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n90,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n89,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n88,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n87,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n86,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n82,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n73,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n72,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n68,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n56,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n55,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n54,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n52,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n51,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n50,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n48,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n46,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n44,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n36,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n28,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n20,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n18,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n10,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n8,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n6,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n4,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n3,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n883,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n139,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n138,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n137,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n11, alu_adder_out_57_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n160,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n950,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n988,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n750,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n749,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n748,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n605, alu_adder_out_22_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n889,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n891,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n494,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n32, alu_adder_out_36_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n294,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n293,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n275,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n274,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n273,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n19, alu_adder_out_49_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n241,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n240,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n239,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n17, alu_adder_out_51_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n411,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n410,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n409,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n27, alu_adder_out_41_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n462,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n460,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n30, alu_adder_out_38_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n394,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n393,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n392,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n26, alu_adder_out_42_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n377,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n376,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n375,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n25, alu_adder_out_43_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n633,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n840,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n927,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n962,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n530,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n529,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n528,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n34, alu_adder_out_34_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n513,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n512,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n511,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n33, alu_adder_out_35_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n497,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n479,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n478,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n477,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n31, alu_adder_out_37_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n207,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n206,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n205,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n15, alu_adder_out_53_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n343,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n342,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n341,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n23, alu_adder_out_45_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n326,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n325,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n324,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n22, alu_adder_out_46_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n767,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n908,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n635,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n737,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n778,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n914,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n932,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n634,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n736,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n790,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n814,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n994,
         alu_addsub_rs2_data_6_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n224,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n223,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n222,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n16, alu_adder_out_52_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n9,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n124,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n105,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n103,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n641,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n639,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n825,
         alu_addsub_rs2_data_15_,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n838,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n846,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n844,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n841,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n960,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n945,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n931,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n929,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n928,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n975,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n969,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n964,
         alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n963,
         alu_addsub_rs2_data_1_, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579;
  wire   [0:62] alu_adder_out;
  wire   [0:63] alu_addsub_rs2_data;

  HDEXNOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U974 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n915), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n619), .Z(alu_adder_out[8])
         );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U989 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n926), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n916), .B(n1864), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n915) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U988 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n926), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n620), .Z(alu_adder_out[7])
         );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U695 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n983), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n682), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n600) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U727 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n985), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n708), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n602) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U928 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n998), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n870), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n615) );
  HDEXNOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U932 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n882), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n616), .Z(alu_adder_out[11]) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U743 ( .A1(n2167), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n721), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n603) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U102 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n569), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n107), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n10) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U62 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n82), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n73), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n8) );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U237 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n268), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n233), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n234), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n228) );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U397 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n369), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n404), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n370), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n364) );
  HDNOR2D2 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U464 ( .A1(n2120), .A2(
        byp_alu_rs1_data_e[40]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n412) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U747 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n735), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n604), .Z(alu_adder_out[23]) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U942 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n999), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n881), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n616) );
  HDEXNOR2DL alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U1037 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n961), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n624), .Z(alu_adder_out[3])
         );
  HDNAN2DL alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U920 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n885), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n863), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n861) );
  HDNAN2DL alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U302 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n579), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n277), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n20) );
  HDNOR2D2 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U264 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_18_), .A2(
        byp_alu_rs1_data_e[50]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n242) );
  HDNAN2D2 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U643 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n662), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n640), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n638) );
  HDNOR2D2 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U898 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n854), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n847), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n845) );
  HDNOR2D2 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U902 ( .A1(
        alu_addsub_rs2_data[14]), .A2(byp_alu_rs1_data_e[14]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n847) );
  HDNOR2D2 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U236 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n267), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n233), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n227) );
  HDNOR2D2 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U316 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n331), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n301), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n299) );
  HDNOR2D2 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U384 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_12_), .A2(
        byp_alu_rs1_data_e[44]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n344) );
  HDNOR2D2 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U476 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n437), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n471), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n435) );
  HDNOR2D2 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U761 ( .A1(n2111), .A2(
        byp_alu_rs1_data_e[23]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n725) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U779 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n761), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n606), .Z(alu_adder_out[21]) );
  HDEXNOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U960 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n904), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n618), .Z(alu_adder_out[9])
         );
  HDEXNOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U946 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n893), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n617), .Z(alu_adder_out[10]) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U683 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n683), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n600), .Z(alu_adder_out[27]) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U715 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n709), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n602), .Z(alu_adder_out[25]) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U859 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n826), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n611), .Z(alu_adder_out[16]) );
  HDEXNOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U904 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n860), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n614), .Z(alu_adder_out[13]) );
  HDEXNOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U918 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n871), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n615), .Z(alu_adder_out[12]) );
  HDEXNOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U891 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n849), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n613), .Z(alu_adder_out[14]) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U827 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n800), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n609), .Z(alu_adder_out[18]) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U731 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n722), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n603), .Z(alu_adder_out[24]) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U651 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n657), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n598), .Z(alu_adder_out[29]) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U637 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n644), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n597), .Z(alu_adder_out[30]) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U699 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n696), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n601), .Z(alu_adder_out[26]) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U667 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n670), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n599), .Z(alu_adder_out[28]) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U795 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n774), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n607), .Z(alu_adder_out[20]) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U811 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n787), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n608), .Z(alu_adder_out[19]) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U10 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n52), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n6), .Z(alu_adder_out[62])
         );
  HDNOR2D2 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U396 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n403), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n369), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n363) );
  HDNOR2D2 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U556 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n531), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n505), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n499) );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U975 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n926), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n905), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n906), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n904) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U956 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n1000), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n892), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n617) );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U961 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n926), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n894), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n895), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n893) );
  HDNOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U733 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n738), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n712), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n710) );
  HDAOI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U876 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n839), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n995), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n828), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n826) );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U919 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n926), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n861), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n862), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n860) );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U933 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n926), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n872), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n873), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n871) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U934 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n885), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n999), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n872) );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U905 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n926), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n850), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n851), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n849) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U906 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n852), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n885), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n850) );
  HDAOI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U844 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n839), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n801), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n802), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n800) );
  HDAOI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U748 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n839), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n723), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n724), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n722) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U663 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n981), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n652), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n598) );
  HDAOI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U668 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n839), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n658), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n659), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n657) );
  HDNOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U669 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n738), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n660), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n658) );
  HDAOI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U652 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n839), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n645), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n646), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n644) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U655 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n649), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n688), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n647) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U711 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n984), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n695), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n601) );
  HDAOI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U716 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n839), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n697), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n698), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n696) );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U718 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n739), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n699), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n700), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n698) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U679 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n982), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n669), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n599) );
  HDAOI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U684 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n839), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n671), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n672), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n670) );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U686 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n739), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n673), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n674), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n672) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U687 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n688), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n983), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n673) );
  HDAOI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U812 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n839), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n775), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n776), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n774) );
  HDAOI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U828 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n839), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n792), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n793), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n787) );
  HDAOI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U351 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n432), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n329), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n330), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n328) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U350 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n329), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n431), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n327) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U246 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n256), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n18), .Z(alu_adder_out[50])
         );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U430 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n431), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n397), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n395) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U270 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n4), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n261), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n259) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U86 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n120), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n10), .Z(alu_adder_out[58])
         );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U446 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n426), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n28), .Z(alu_adder_out[40])
         );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U45 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_29_), .A2(
        byp_alu_rs1_data_e[61]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n68) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U46 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n86), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n8), .Z(alu_adder_out[60])
         );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U190 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n4), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n193), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n191) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U125 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_25_), .A2(
        byp_alu_rs1_data_e[57]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n136) );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U157 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n196), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n165), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n166), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n164) );
  HDAOI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U159 ( .A1(n2487), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n185), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n168), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n166) );
  HDAOI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U199 ( .A1(n2488), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n219), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n202), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n196) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U205 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_21_), .A2(
        byp_alu_rs1_data_e[53]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n204) );
  HDAOI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U239 ( .A1(n2495), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n253), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n236), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n234) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U245 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_19_), .A2(
        byp_alu_rs1_data_e[51]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n238) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U285 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_17_), .A2(
        byp_alu_rs1_data_e[49]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n272) );
  HDAOI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U319 ( .A1(n2489), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n321), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n304), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n302) );
  HDAOI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U359 ( .A1(n2493), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n355), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n338), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n332) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U365 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_13_), .A2(
        byp_alu_rs1_data_e[45]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n340) );
  HDAOI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U399 ( .A1(n2490), .A2(
        n2194), .B(n2125), .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n370)
         );
  HDAOI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U519 ( .A1(n2494), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n491), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n474), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n472) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U150 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n4), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n159), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n157) );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U678 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n668), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n682), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n669), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n663) );
  HDNOR2D2 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U926 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n869), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n880), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n863) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U106 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n137), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n11), .Z(alu_adder_out_57_)
         );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U122 ( .A1(n2484), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n136), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n11) );
  HDNOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U128 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n157), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n140), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n138) );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U129 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n158), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n140), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n141), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n139) );
  HDNOR2D2 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U930 ( .A1(n2168), .A2(
        byp_alu_rs1_data_e[12]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n869) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U763 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n748), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n605), .Z(alu_adder_out_22_) );
  HDAOI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U780 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n839), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n749), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n750), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n748) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U775 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n988), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n747), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n605) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U526 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n494), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n32), .Z(alu_adder_out_36_)
         );
  HDNAN2DL alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U542 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n591), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n481), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n32) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U266 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n273), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n19), .Z(alu_adder_out_49_)
         );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U282 ( .A1(n2485), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n272), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n19) );
  HDNOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U288 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n293), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n276), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n274) );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U289 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n294), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n276), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n277), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n275) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U226 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n239), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n17), .Z(alu_adder_out_51_)
         );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U242 ( .A1(n2495), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n238), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n17) );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U249 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n260), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n242), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n243), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n241) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U426 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n409), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n27), .Z(alu_adder_out_41_)
         );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U442 ( .A1(n2486), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n408), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n27) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U486 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n460), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n30), .Z(alu_adder_out_38_)
         );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U406 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n392), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n26), .Z(alu_adder_out_42_)
         );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U386 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n375), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n25), .Z(alu_adder_out_43_)
         );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U409 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n396), .A2(n1790), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n379), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n377) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U566 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n528), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n34), .Z(alu_adder_out_34_)
         );
  HDNAN2DL alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U582 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n593), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n515), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n34) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U546 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n511), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n33), .Z(alu_adder_out_35_)
         );
  HDNAN2DL alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U562 ( .A1(n1770), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n510), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n33) );
  HDNOR2DL alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U568 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n531), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n514), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n512) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U506 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n477), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n31), .Z(alu_adder_out_37_)
         );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U522 ( .A1(n2494), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n476), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n31) );
  HDNOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U528 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n497), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n480), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n478) );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U529 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n498), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n480), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n481), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n479) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U186 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n205), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n15), .Z(alu_adder_out_53_)
         );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U202 ( .A1(n2488), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n204), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n15) );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U209 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n226), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n208), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n209), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n207) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U346 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n341), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n23), .Z(alu_adder_out_45_)
         );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U362 ( .A1(n2493), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n340), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n23) );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U369 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n362), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n344), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n345), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n343) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U326 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n324), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n22), .Z(alu_adder_out_46_)
         );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U342 ( .A1(n1791), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n311), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n22) );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U806 ( .A1(n1748), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n778), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n773), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n767) );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U638 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n840), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n634), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n635), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n633) );
  HDNOR2DL alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U813 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n790), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n777), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n775) );
  HDEXOR2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U206 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n222), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n16), .Z(alu_adder_out_52_)
         );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U222 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n575), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n209), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n16) );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U89 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n124), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n106), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n107), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n105) );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U646 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n642), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n652), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n643), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n641) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U230 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n4), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n227), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n225) );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U899 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n847), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n855), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n848), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n846) );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U1032 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n950), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n960), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n951), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n945) );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U1008 ( .A1(n2108), 
        .A2(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n938), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n933), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n931) );
  HDOAI21D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U1053 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n969), .A2(n1736), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n966), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n964) );
  HDNOR2D2 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U889 ( .A1(n2146), .A2(
        byp_alu_rs1_data_e[15]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n837) );
  HDNAN2D2 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U931 ( .A1(
        alu_addsub_rs2_data[12]), .A2(byp_alu_rs1_data_e[12]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n870) );
  HDNAN2D2 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U636 ( .A1(
        alu_addsub_rs2_data[31]), .A2(byp_alu_rs1_data_e[31]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n632) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U262 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n577), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n243), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n18) );
  HDNAN2DL alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U633 ( .A1(n2496), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n632), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n596) );
  HDNAN2D2 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U38 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n82), .A2(n2482), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n55) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U719 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n714), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n985), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n699) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U22 ( .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n565), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n51), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n6) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U25 ( .A1(
        alu_addsub_rs2_data[62]), .A2(byp_alu_rs1_data_e[62]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n51) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U82 ( .A1(n2483), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n102), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n9) );
  HDNAN2D1 alu_addsub_adder_add_24_2_DP_OP_282_4997_7_U422 ( .A1(n1869), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n379), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n26) );
  HDNAN2D1 U1562 ( .A1(n2700), .A2(byp_alu_rs1_data_e[16]), .Z(n2996) );
  HDNAN2D1 U1563 ( .A1(n2701), .A2(byp_alu_rs1_data_e[17]), .Z(n3005) );
  HDOAI21M20D1 U1564 ( .A1(byp_alu_rs1_data_e[51]), .A2(n2745), .B(n2676), .Z(
        n3311) );
  HDINVD1 U1565 ( .A(n3418), .Z(n3261) );
  HDINVD1 U1566 ( .A(n3445), .Z(n3305) );
  HDOR2D1 U1567 ( .A1(n1744), .A2(n2586), .Z(n2507) );
  HDINVD1 U1568 ( .A(n3474), .Z(n3331) );
  HDNAN2D1 U1569 ( .A1(n2668), .A2(byp_alu_rs1_data_e[23]), .Z(n3339) );
  HDNAN2D1 U1570 ( .A1(n2203), .A2(byp_alu_rs1_data_e[46]), .Z(n3403) );
  HDNOR2D1 U1571 ( .A1(n2506), .A2(n3567), .Z(n3413) );
  HDINVD1 U1572 ( .A(n3458), .Z(n3316) );
  HDINVD1 U1573 ( .A(n3483), .Z(n3340) );
  HDINVD2 U1574 ( .A(n3529), .Z(n3383) );
  HDINVD1 U1575 ( .A(n3535), .Z(n3394) );
  HDAOI211D2 U1576 ( .A1(ecl_shft_shift4_e[2]), .A2(n3354), .B(n3286), .C(
        n3285), .Z(n3310) );
  HDOAI211D2 U1577 ( .A1(n3340), .A2(n2655), .B(n2021), .C(n3339), .Z(n3449)
         );
  HDNAN2D1 U1578 ( .A1(n2700), .A2(byp_alu_rs1_data_e[39]), .Z(n2021) );
  HDOA211D2 U1579 ( .A1(n3513), .A2(n2655), .B(n3363), .C(n3362), .Z(n3478) );
  HDOR2D1 U1580 ( .A1(ecl_shft_enshift_e_l), .A2(byp_alu_rs2_data_e[4]), .Z(
        n2199) );
  HDINVD4 U1581 ( .A(byp_alu_rs2_data_e[5]), .Z(n1820) );
  HDNAN2D4 U1582 ( .A1(n2712), .A2(ecl_shft_op32_e), .Z(n2659) );
  HDNAN2D1 U1583 ( .A1(n2701), .A2(byp_alu_rs1_data_e[25]), .Z(n3123) );
  HDINVD1 U1584 ( .A(n3311), .Z(n3062) );
  HDNAN2D1 U1585 ( .A1(n2700), .A2(byp_alu_rs1_data_e[29]), .Z(n3201) );
  HDNOR2D1 U1586 ( .A1(n2741), .A2(ecl_shft_enshift_e_l), .Z(n3535) );
  HDINVD1 U1587 ( .A(byp_alu_rs1_data_e[13]), .Z(n2741) );
  HDINVD1 U1588 ( .A(n1768), .Z(n2698) );
  HDINVD1 U1589 ( .A(byp_alu_rs1_data_e[4]), .Z(n2235) );
  HDNAN2D1 U1590 ( .A1(n2203), .A2(byp_alu_rs1_data_e[22]), .Z(n3085) );
  HDNAN2D1 U1591 ( .A1(n2699), .A2(byp_alu_rs1_data_e[26]), .Z(n3142) );
  HDINVD1 U1592 ( .A(byp_alu_rs1_data_e[6]), .Z(n2717) );
  HDNAN2D4 U1593 ( .A1(n2684), .A2(ecl_shft_shift4_e[1]), .Z(n3040) );
  HDOA21D1 U1594 ( .A1(n2119), .A2(n3422), .B(n2996), .Z(n3184) );
  HDAND2D1 U1595 ( .A1(alu_addsub_rs2_data[32]), .A2(byp_alu_rs1_data_e[32]), 
        .Z(n2469) );
  HDNOR2D1 U1596 ( .A1(n2136), .A2(byp_alu_rs1_data_e[32]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n560) );
  HDINVD1 U1597 ( .A(n3367), .Z(n3219) );
  HDAOI21D1 U1598 ( .A1(n1770), .A2(n2156), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n508), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n506) );
  HDOAI21M20D1 U1599 ( .A1(n3108), .A2(n2681), .B(n3107), .Z(n3317) );
  HDEXOR2DL U1600 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[39]), .Z(
        n2182) );
  HDOR2D1 U1601 ( .A1(n3361), .A2(n2702), .Z(n2084) );
  HDAOI211D2 U1602 ( .A1(n1782), .A2(n3177), .B(n3176), .C(n2016), .Z(n3345)
         );
  HDNOR2D1 U1603 ( .A1(n3175), .A2(n1773), .Z(n2016) );
  HDINVD1 U1604 ( .A(n3389), .Z(n3198) );
  HDAOI211D2 U1605 ( .A1(n3461), .A2(ecl_shft_shift4_e[1]), .B(n3386), .C(
        n3385), .Z(n1779) );
  HDAND4D1 U1606 ( .A1(n2448), .A2(n2449), .A3(n1774), .A4(n2450), .Z(n3406)
         );
  HDNOR2D1 U1607 ( .A1(n2001), .A2(n2706), .Z(n1962) );
  HDINVD1 U1608 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n243), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n253) );
  HDOR2D1 U1609 ( .A1(n3490), .A2(n3533), .Z(n2036) );
  HDAOI211D2 U1610 ( .A1(ecl_shft_shift4_e[0]), .A2(n3543), .B(n3507), .C(
        n3506), .Z(n3525) );
  HDNOR2D1 U1611 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n161), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n93), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n91) );
  HDEXOR2D1 U1612 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[61]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_29_) );
  HDINVD1 U1613 ( .A(ecl_shft_shift1_e[0]), .Z(n2751) );
  HDOR2D1 U1614 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_29_), .A2(
        byp_alu_rs1_data_e[61]), .Z(n2482) );
  HDNAN2D1 U1615 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n569), .A2(
        n2483), .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n97) );
  HDOA21M20D2 U1616 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n364), 
        .A2(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n299), .B(n2133), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n298) );
  HDNAN2D2 U1617 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n227), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n163), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n161) );
  HDNAN2D1 U1618 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n95), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n48), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n46) );
  HDINVD1 U1619 ( .A(n2807), .Z(n2767) );
  HDOR2D1 U1620 ( .A1(n2977), .A2(n3431), .Z(n2807) );
  HDOA211D1 U1621 ( .A1(n2892), .A2(n2704), .B(n2835), .C(n2834), .Z(n2881) );
  HDINVD1 U1622 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n560), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n595) );
  HDINVD1 U1623 ( .A(byp_alu_rs1_data_e[34]), .Z(n3438) );
  HDOA22D1 U1624 ( .A1(n3334), .A2(n3561), .B1(n3333), .B2(n1789), .Z(n2249)
         );
  HDNOR2D1 U1625 ( .A1(n3341), .A2(n2708), .Z(n3306) );
  HDOA222D1 U1626 ( .A1(n3343), .A2(n3560), .B1(n3334), .B2(n3576), .C1(n3325), 
        .C2(n2686), .Z(n2073) );
  HDINVD1 U1627 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n429), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n431) );
  HDINVD1 U1628 ( .A(byp_alu_rs1_data_e[40]), .Z(n3346) );
  HDAOI211D2 U1629 ( .A1(ecl_shft_shift4_e[3]), .A2(n2508), .B(n3442), .C(
        n3441), .Z(n3468) );
  HDNOR2D1 U1630 ( .A1(n3487), .A2(n2456), .Z(n2513) );
  HDNAN2D1 U1631 ( .A1(n1792), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n175), .Z(n2233) );
  HDNOR2D1 U1632 ( .A1(n3500), .A2(n3563), .Z(n2034) );
  HDNAN2D1 U1633 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n170), .A2(
        n2487), .Z(n2313) );
  HDOR2D1 U1634 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_25_), .A2(
        byp_alu_rs1_data_e[57]), .Z(n2484) );
  HDEXOR2D1 U1635 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[57]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_25_) );
  HDAOI211D2 U1636 ( .A1(ecl_shft_shift4_e[0]), .A2(n3570), .B(n3488), .C(
        n3489), .Z(n3508) );
  HDNOR2D1 U1637 ( .A1(n3487), .A2(n2704), .Z(n3488) );
  HDEXOR2D1 U1638 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[58]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_26_) );
  HDNAN2D1 U1639 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_26_), 
        .A2(byp_alu_rs1_data_e[58]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n107) );
  HDNAN2D1 U1640 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_27_), 
        .A2(byp_alu_rs1_data_e[59]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n102) );
  HDNAN2D1 U1641 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_28_), 
        .A2(byp_alu_rs1_data_e[60]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n73) );
  HDINVD2 U1642 ( .A(n3548), .Z(n3574) );
  HDNOR2D1 U1643 ( .A1(n2751), .A2(ecl_shft_lshift_e_l), .Z(n2688) );
  HDOA21M10DL U1644 ( .A2(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n73), 
        .A1(n2482), .B(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n68), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n56) );
  HDNOR2D1 U1645 ( .A1(alu_addsub_rs2_data[62]), .A2(byp_alu_rs1_data_e[62]), 
        .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n50) );
  HDNOR2D1 U1646 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n46), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n162), .Z(n2270) );
  HDNOR2D1 U1647 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n55), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n50), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n48) );
  HDNOR2D1 U1648 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n161), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n46), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n44) );
  HDEXOR2D1 U1649 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[62]), .Z(
        alu_addsub_rs2_data[62]) );
  HDINVBD4 U1650 ( .A(byp_alu_rs2_data_e[16]), .Z(n1983) );
  HDINVD12 U1651 ( .A(ifu_exu_invert_d), .Z(n1747) );
  HDNAN2D1 U1652 ( .A1(n2110), .A2(byp_alu_rs1_data_e[23]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n726) );
  HDNOR2D1 U1653 ( .A1(alu_addsub_rs2_data[8]), .A2(byp_alu_rs1_data_e[8]), 
        .Z(n1892) );
  HDEXOR2D1 U1654 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[8]), .Z(
        alu_addsub_rs2_data[8]) );
  HDNAN2D1 U1655 ( .A1(n2743), .A2(byp_alu_rs1_data_e[18]), .Z(n3437) );
  HDINVD1 U1656 ( .A(n2822), .Z(n2715) );
  HDINVBD2 U1657 ( .A(byp_alu_rs2_data_e[15]), .Z(n1816) );
  HDINVD1 U1658 ( .A(n3437), .Z(n2786) );
  HDINVD1 U1659 ( .A(byp_alu_rs1_data_e[18]), .Z(n1811) );
  HDINVD2 U1660 ( .A(byp_alu_rs2_data_e[18]), .Z(n1874) );
  HDNOR2D1 U1661 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n651), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n642), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n640) );
  HDOAI21M20D1 U1662 ( .A1(byp_alu_rs1_data_e[33]), .A2(n2745), .B(n2659), .Z(
        n3019) );
  HDNAN2D1 U1663 ( .A1(n2700), .A2(byp_alu_rs1_data_e[20]), .Z(n3059) );
  HDNAN2D1 U1664 ( .A1(n2203), .A2(byp_alu_rs1_data_e[23]), .Z(n3095) );
  HDEXOR2DL U1665 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[39]), .Z(
        n2183) );
  HDINVD1 U1666 ( .A(ecl_shft_shift4_e[0]), .Z(n1750) );
  HDINVD1 U1667 ( .A(n2710), .Z(n1751) );
  HDNAN2D1 U1668 ( .A1(n2203), .A2(byp_alu_rs1_data_e[37]), .Z(n2511) );
  HDINVD1 U1669 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n238), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n236) );
  HDNAN2D1 U1670 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n579), .A2(
        n2485), .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n267) );
  HDINVD1 U1671 ( .A(ecl_shft_shift4_e[3]), .Z(n1749) );
  HDINVD1 U1672 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n175), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n185) );
  HDINVD1 U1673 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n170), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n168) );
  HDINVD1 U1674 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n306), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n304) );
  HDNAN2D1 U1675 ( .A1(n2818), .A2(ecl_shft_shift4_e[2]), .Z(n2736) );
  HDINVBD4 U1676 ( .A(ifu_exu_invert_d), .Z(n1746) );
  HDINVD1 U1677 ( .A(byp_alu_rs1_data_e[2]), .Z(n1796) );
  HDNOR2D1 U1678 ( .A1(n2000), .A2(byp_alu_rs1_data_e[4]), .Z(n2464) );
  HDOA211D1 U1679 ( .A1(n3340), .A2(n2685), .B(n2730), .C(n3339), .Z(n2804) );
  HDEXOR2D1 U1680 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[7]), .Z(
        alu_addsub_rs2_data[7]) );
  HDEXOR2DL U1681 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[9]), .Z(
        n1999) );
  HDINVD1 U1682 ( .A(n3521), .Z(n2907) );
  HDAND2D1 U1683 ( .A1(n2729), .A2(n2728), .Z(n2928) );
  HDINVD1 U1684 ( .A(n3498), .Z(n3108) );
  HDINVD1 U1685 ( .A(n3422), .Z(n2866) );
  HDINVD1 U1686 ( .A(n3505), .Z(n3124) );
  HDINVD1 U1687 ( .A(n3513), .Z(n3143) );
  HDINVD1 U1688 ( .A(n3436), .Z(n2888) );
  HDAOI211D1 U1689 ( .A1(n2959), .A2(n3458), .B(n2926), .C(n2925), .Z(n2983)
         );
  HDINVD1 U1690 ( .A(ecl_shft_shift1_e[1]), .Z(n2765) );
  HDINVD1 U1691 ( .A(n3464), .Z(n3320) );
  HDINVD1 U1692 ( .A(n1882), .Z(n1883) );
  HDINVD1 U1693 ( .A(n3314), .Z(n3178) );
  HDAND2D1 U1694 ( .A1(alu_addsub_rs2_data[34]), .A2(byp_alu_rs1_data_e[34]), 
        .Z(n2156) );
  HDOR2D1 U1695 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_7_), .A2(
        byp_alu_rs1_data_e[39]), .Z(n2492) );
  HDNAN2D1 U1696 ( .A1(n2183), .A2(byp_alu_rs1_data_e[39]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n442) );
  HDINVD1 U1697 ( .A(n2447), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n423) );
  HDINVD1 U1698 ( .A(n1807), .Z(n2588) );
  HDNOR2D1 U1699 ( .A1(n2583), .A2(n3288), .Z(n2585) );
  HDNOR2D1 U1700 ( .A1(n2358), .A2(n2364), .Z(n1914) );
  HDINVD1 U1701 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n340), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n338) );
  HDINVD1 U1702 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n345), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n355) );
  HDNAN2D1 U1703 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_15_), 
        .A2(byp_alu_rs1_data_e[47]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n306) );
  HDAOI211D2 U1704 ( .A1(ecl_shft_shift4_e[1]), .A2(n3457), .B(n3420), .C(
        n3419), .Z(n3451) );
  HDINVD1 U1705 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n267), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n261) );
  HDNOR2D1 U1706 ( .A1(n3575), .A2(n2710), .Z(n3456) );
  HDNAN2D1 U1707 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_23_), 
        .A2(byp_alu_rs1_data_e[55]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n170) );
  HDOR2D1 U1708 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_23_), .A2(
        byp_alu_rs1_data_e[55]), .Z(n2487) );
  HDINVD2 U1709 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n174), .Z(
        n1792) );
  HDINVD1 U1710 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n141), .Z(
        n1784) );
  HDINVD2 U1711 ( .A(n2121), .Z(n2005) );
  HDINVD1 U1712 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n161), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n159) );
  HDNAN2D1 U1713 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n571), .A2(
        n2484), .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n127) );
  HDOA211D1 U1714 ( .A1(n3383), .A2(n2299), .B(n3382), .C(n3381), .Z(n2123) );
  HDAND2D1 U1715 ( .A1(n3466), .A2(n3465), .Z(n3540) );
  HDINVD1 U1716 ( .A(n3556), .Z(n3515) );
  HDOA211D1 U1717 ( .A1(n3553), .A2(n2694), .B(n3403), .C(n1730), .Z(n1877) );
  HDNAN2D1 U1718 ( .A1(n2698), .A2(byp_alu_rs1_data_e[59]), .Z(n2545) );
  HDAOI22D1 U1719 ( .A1(n3536), .A2(n3445), .B1(n2138), .B2(
        byp_alu_rs1_data_e[51]), .Z(n3446) );
  HDAOI211D2 U1720 ( .A1(n2138), .A2(byp_alu_rs1_data_e[47]), .B(n3413), .C(
        n3412), .Z(n3524) );
  HDNOR2D1 U1721 ( .A1(n2299), .A2(n3565), .Z(n3412) );
  HDINVD1 U1722 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n56), .Z(n1752) );
  HDOR2D1 U1723 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n89), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n55), .Z(n2150) );
  HDINVD2 U1724 ( .A(ecl_shft_lshift_e_l), .Z(n3578) );
  HDINVD1 U1725 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n976), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n1010) );
  HDNAN2D1 U1726 ( .A1(byp_alu_rs1_data_e[0]), .A2(ecl_alu_cin_e), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n977) );
  HDOA211D1 U1727 ( .A1(n2887), .A2(n2704), .B(n2821), .C(n2820), .Z(n2455) );
  HDOA211D1 U1728 ( .A1(n2887), .A2(n2704), .B(n2821), .C(n2820), .Z(n2864) );
  HDINVD2 U1729 ( .A(byp_alu_rs2_data_e[13]), .Z(n2164) );
  HDOA211D1 U1730 ( .A1(n2892), .A2(n2456), .B(n2891), .C(n2890), .Z(n2941) );
  HDNAN2D1 U1731 ( .A1(n2174), .A2(byp_alu_rs1_data_e[14]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n848) );
  HDBUFD1 U1732 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n838), .Z(
        n2177) );
  HDNOR3D2 U1733 ( .A1(n2204), .A2(n2980), .A3(n2181), .Z(n3158) );
  HDNOR2D1 U1734 ( .A1(n2765), .A2(n3578), .Z(n3549) );
  HDOA211D1 U1735 ( .A1(n3137), .A2(n2710), .B(n2964), .C(n2963), .Z(n3012) );
  HDNOR2D1 U1736 ( .A1(n2998), .A2(n2997), .Z(n3038) );
  HDOA211D1 U1737 ( .A1(n3137), .A2(n2706), .B(n3024), .C(n3023), .Z(n3075) );
  HDNOR2D1 U1738 ( .A1(n3042), .A2(n3041), .Z(n3094) );
  HDAO21M10DL U1739 ( .A2(n2315), .A1(n2185), .B(n2316), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n750) );
  HDNOR2D1 U1740 ( .A1(n3079), .A2(n3078), .Z(n3106) );
  HDAOI211D2 U1741 ( .A1(ecl_shft_shift4_e[0]), .A2(n3092), .B(n3091), .C(
        n3090), .Z(n3117) );
  HDNOR2D1 U1742 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n738), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n699), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n697) );
  HDNOR2D1 U1743 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n738), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n673), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n671) );
  HDNOR2D1 U1744 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n738), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n647), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n645) );
  HDNAN2D1 U1745 ( .A1(n1978), .A2(byp_alu_rs1_data_e[30]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n643) );
  HDNOR2D1 U1746 ( .A1(n3257), .A2(n2456), .Z(n3263) );
  HDEXOR2DL U1747 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[33]), .Z(
        n2151) );
  HDINVD1 U1748 ( .A(n2156), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n515) );
  HDOR2D1 U1749 ( .A1(n2141), .A2(byp_alu_rs1_data_e[35]), .Z(n1770) );
  HDOA211D1 U1750 ( .A1(n2706), .A2(n3219), .B(n2003), .C(n2004), .Z(n3324) );
  HDNOR2D1 U1751 ( .A1(n3332), .A2(n2705), .Z(n2328) );
  HDINVD1 U1752 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n480), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n591) );
  HDOA22D1 U1753 ( .A1(n3334), .A2(n3560), .B1(n3333), .B2(n3563), .Z(n1931)
         );
  HDEXOR2DL U1754 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[37]), .Z(
        n1934) );
  HDNAN2D1 U1755 ( .A1(n1967), .A2(byp_alu_rs1_data_e[37]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n476) );
  HDOR2D1 U1756 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_5_), .A2(
        byp_alu_rs1_data_e[37]), .Z(n2494) );
  HDOAI22M10D1 U1757 ( .A1(n2503), .A2(n3343), .B1(n2686), .B2(n3342), .Z(
        n2581) );
  HDOR2D1 U1758 ( .A1(n3388), .A2(n3561), .Z(n2083) );
  HDEXOR2DL U1759 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[41]), .Z(
        n2186) );
  HDOA22D1 U1760 ( .A1(n3369), .A2(n2702), .B1(n3388), .B2(n3560), .Z(n2056)
         );
  HDINVD1 U1761 ( .A(n2194), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n379) );
  HDOR2D1 U1762 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_11_), .A2(
        byp_alu_rs1_data_e[43]), .Z(n2490) );
  HDNOR2D1 U1763 ( .A1(n2359), .A2(n1783), .Z(n2411) );
  HDEXOR2DL U1764 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[44]), .Z(
        n1980) );
  HDINVD1 U1765 ( .A(n2689), .Z(n1764) );
  HDINVD1 U1766 ( .A(n1783), .Z(n1745) );
  HDINVD1 U1767 ( .A(n2689), .Z(n1765) );
  HDEXOR2DL U1768 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[46]), .Z(
        n1904) );
  HDINVD1 U1769 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n310), .Z(
        n1791) );
  HDNAN2D1 U1770 ( .A1(n2104), .A2(byp_alu_rs1_data_e[46]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n311) );
  HDINVD1 U1771 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n276), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n579) );
  HDAOI211D2 U1772 ( .A1(ecl_shft_shift4_e[2]), .A2(n2508), .B(n3405), .C(
        n3404), .Z(n3427) );
  HDINVD1 U1773 ( .A(byp_alu_rs1_data_e[48]), .Z(n3414) );
  HDEXOR2DL U1774 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[50]), .Z(
        n1861) );
  HDINVD1 U1775 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n242), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n577) );
  HDNAN2D1 U1776 ( .A1(n1862), .A2(byp_alu_rs1_data_e[50]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n243) );
  HDINVD1 U1777 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n208), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n575) );
  HDEXOR2DL U1778 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[52]), .Z(
        n1808) );
  HDOA22D1 U1779 ( .A1(n3491), .A2(n3560), .B1(n3490), .B2(n3563), .Z(n1921)
         );
  HDOA22D1 U1780 ( .A1(n3469), .A2(n2702), .B1(n3468), .B2(n3533), .Z(n1920)
         );
  HDINVD1 U1781 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n209), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n219) );
  HDINVD1 U1782 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n204), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n202) );
  HDEXOR2D1 U1783 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[56]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_24_) );
  HDAOI211D2 U1784 ( .A1(n3556), .A2(ecl_shft_shift4_e[0]), .B(n3480), .C(
        n3479), .Z(n3500) );
  HDNOR2D1 U1785 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n161), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n127), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n125) );
  HDNOR2D1 U1786 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_26_), 
        .A2(byp_alu_rs1_data_e[58]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n106) );
  HDOR2D1 U1787 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_27_), .A2(
        byp_alu_rs1_data_e[59]), .Z(n2483) );
  HDEXOR2D1 U1788 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[59]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_27_) );
  HDINVD1 U1789 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n96), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n94) );
  HDEXOR2D1 U1790 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[60]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_28_) );
  HDNOR2D1 U1791 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_28_), 
        .A2(byp_alu_rs1_data_e[60]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n72) );
  HDAO211DL U1792 ( .A1(n2284), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_29_), .B(n2285), .C(
        n2286), .Z(n2297) );
  HDINVD1 U1793 ( .A(ecl_alu_log_sel_and_e), .Z(n2757) );
  HDNOR2D4 U1794 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n429), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n297), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n4) );
  HDEXOR2DL U1795 ( .A1(byp_alu_rs2_data_e[63]), .A2(ifu_exu_invert_d), .Z(
        alu_addsub_rs2_data[63]) );
  HDINVD8 U1796 ( .A(n1772), .Z(n2703) );
  HDEXOR2DL U1797 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[1]), .Z(
        n2176) );
  HDINVD1 U1798 ( .A(n2688), .Z(n1726) );
  HDINVD1 U1799 ( .A(n2767), .Z(n1727) );
  HDEXOR2DL U1800 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[2]), .Z(
        n2394) );
  HDEXOR2DL U1801 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[3]), .Z(
        n2334) );
  HDEXOR2D1 U1802 ( .A1(byp_alu_rs2_data_e[4]), .A2(ifu_exu_invert_d), .Z(
        n2000) );
  HDEXOR2DL U1803 ( .A1(ifu_exu_invert_d), .A2(n1742), .Z(n2160) );
  HDEXOR2DL U1804 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[6]), .Z(
        n1880) );
  HDEXOR2DL U1805 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[6]), .Z(
        n2193) );
  HDEXOR2DL U1806 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[7]), .Z(
        n2197) );
  HDEXOR2DL U1807 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[8]), .Z(
        n2189) );
  HDEXOR2DL U1808 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[10]), .Z(
        n2274) );
  HDEXOR2DL U1809 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[11]), .Z(
        n2172) );
  HDEXOR2DL U1810 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[12]), .Z(
        n2169) );
  HDEXOR2DL U1811 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[14]), .Z(
        n2175) );
  HDEXOR2DL U1812 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[15]), .Z(
        n2145) );
  HDOAI21M20DL U1813 ( .A1(n2569), .A2(n1794), .B(n2570), .Z(n2565) );
  HDEXOR2DL U1814 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[18]), .Z(
        n2148) );
  HDEXOR2DL U1815 ( .A1(byp_alu_rs2_data_e[19]), .A2(ifu_exu_invert_d), .Z(
        n1885) );
  HDEXOR2DL U1816 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[20]), .Z(
        n2170) );
  HDEXOR2DL U1817 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[22]), .Z(
        n1804) );
  HDEXOR2DL U1818 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[22]), .Z(
        n2178) );
  HDOA21M20D1 U1819 ( .A1(n2531), .A2(n2110), .B(n2532), .Z(n2537) );
  HDEXOR2DL U1820 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[25]), .Z(
        n2007) );
  HDEXOR2DL U1821 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[26]), .Z(
        n2117) );
  HDEXOR2DL U1822 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[27]), .Z(
        n1867) );
  HDEXOR2DL U1823 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[28]), .Z(
        n1976) );
  HDEXOR2DL U1824 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[29]), .Z(
        n1969) );
  HDEXOR2DL U1825 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[30]), .Z(
        n1979) );
  HDINVBD2 U1826 ( .A(n3278), .Z(n2683) );
  HDEXNOR2D1 U1827 ( .A1(n2012), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n36), .Z(n1759) );
  HDINVD1 U1828 ( .A(n2689), .Z(n1758) );
  HDINVD1 U1829 ( .A(n1785), .Z(n1757) );
  HDEXNOR2DL U1830 ( .A1(n1873), .A2(byp_alu_rs2_data_e[32]), .Z(n2137) );
  HDEXOR2DL U1831 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[34]), .Z(
        n1958) );
  HDINVD1 U1832 ( .A(byp_alu_rs2_data_e[36]), .Z(n1725) );
  HDNOR2D4 U1833 ( .A1(n3333), .A2(n1783), .Z(n2067) );
  HDOA21D1 U1834 ( .A1(n2418), .A2(ecl_alu_out_sel_shift_e_l), .B(n2432), .Z(
        n2417) );
  HDOA211D1 U1835 ( .A1(n2380), .A2(ecl_alu_out_sel_shift_e_l), .B(n2381), .C(
        n2382), .Z(n2379) );
  HDNAN2M1D1 U1836 ( .A1(n2377), .A2(n2383), .Z(n2382) );
  HDOR2D1 U1837 ( .A1(n3470), .A2(n1789), .Z(n2097) );
  HDOR2D1 U1838 ( .A1(n3470), .A2(n3563), .Z(n1860) );
  HDINVD2 U1839 ( .A(n2311), .Z(n2027) );
  HDEXOR2D1 U1840 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[55]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_23_) );
  HDNOR3D1 U1841 ( .A1(n2032), .A2(n2033), .A3(n1775), .Z(n2031) );
  HDNOR2D1 U1842 ( .A1(n3508), .A2(n1789), .Z(n2033) );
  HDOAI21M20D1 U1843 ( .A1(n2481), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n44), .B(n2268), .Z(n2254)
         );
  HDNOR2D1 U1844 ( .A1(n3573), .A2(n1795), .Z(n2259) );
  HDAO22DL U1845 ( .A1(byp_alu_rs2_data_e[0]), .A2(n2683), .B1(
        alu_adder_out[0]), .B2(n1785), .Z(n2674) );
  HDOAI21M20DL U1846 ( .A1(n2544), .A2(n1924), .B(n2538), .Z(
        alu_byp_rd_data_e[9]) );
  HDNOR2D1 U1847 ( .A1(n2579), .A2(n2499), .Z(n2578) );
  HDOA21D1 U1848 ( .A1(n2222), .A2(ecl_alu_out_sel_shift_e_l), .B(n2234), .Z(
        n2221) );
  HDNOR2D1 U1849 ( .A1(n2373), .A2(n2374), .Z(n2372) );
  HDOA211D1 U1850 ( .A1(n2593), .A2(ecl_alu_out_sel_shift_e_l), .B(n2594), .C(
        n2595), .Z(n2592) );
  HDOR2D1 U1851 ( .A1(n2279), .A2(n2280), .Z(n2278) );
  HDINVD1 U1852 ( .A(ecl_shft_extendbit_e), .Z(n1740) );
  HDNOR2M1D1 U1853 ( .A1(n3283), .A2(n3566), .Z(n2735) );
  HDNAN2D1 U1854 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[23]), .Z(
        n1576) );
  HDOAI211D1 U1855 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[23]), .B(
        byp_alu_rs1_data_e[23]), .C(n1576), .Z(n2134) );
  HDOA21M20D1 U1856 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n689), 
        .A2(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n662), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n665), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n661) );
  HDNOR2D1 U1857 ( .A1(n2709), .A2(n2510), .Z(n1577) );
  HDOAI22D1 U1858 ( .A1(n2585), .A2(n2710), .B1(n2589), .B2(n2456), .Z(n1578)
         );
  HDAOI211D2 U1859 ( .A1(ecl_shft_shift4_e[1]), .A2(n3467), .B(n1577), .C(
        n1578), .Z(n2590) );
  HDOAI21M20DL U1860 ( .A1(n2477), .A2(n1805), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n938), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n936) );
  HDNAN2D1 U1861 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[9]), .Z(n1579) );
  HDOAI211D1 U1862 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[9]), .B(
        byp_alu_rs1_data_e[9]), .C(n1579), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n903) );
  HDAOI22D1 U1863 ( .A1(n3011), .A2(ecl_shft_shift4_e[1]), .B1(
        ecl_shft_shift4_e[2]), .B2(n3084), .Z(n1580) );
  HDNAN2M1D1 U1864 ( .A1(n2456), .A2(n2946), .Z(n1581) );
  HDOA211D1 U1865 ( .A1(n3119), .A2(n2710), .B(n1580), .C(n1581), .Z(n2994) );
  HDOAI22D1 U1866 ( .A1(n3241), .A2(n2706), .B1(n3565), .B2(n3165), .Z(n1582)
         );
  HDOAI22D1 U1867 ( .A1(n3341), .A2(n2456), .B1(n3164), .B2(n2704), .Z(n1583)
         );
  HDNOR2D1 U1868 ( .A1(n1582), .A2(n1583), .Z(n3225) );
  HDNOR2M1D1 U1869 ( .A1(n3295), .A2(n3566), .Z(n1584) );
  HDAOI211D1 U1870 ( .A1(n1786), .A2(n3019), .B(n3288), .C(n1584), .Z(n2748)
         );
  HDNAN2D1 U1871 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[2]), .Z(n1585) );
  HDOAI211D1 U1872 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[2]), .B(
        byp_alu_rs1_data_e[2]), .C(n1585), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n966) );
  HDNOR2M1D1 U1873 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n863), 
        .A2(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n854), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n852) );
  HDNAN2D1 U1874 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[27]), .Z(
        n1586) );
  HDOAI211D1 U1875 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[27]), .B(
        byp_alu_rs1_data_e[27]), .C(n1586), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n682) );
  HDNAN2D1 U1876 ( .A1(n3061), .A2(n1782), .Z(n1587) );
  HDOA211D1 U1877 ( .A1(n3062), .A2(n1773), .B(n3260), .C(n1587), .Z(n3257) );
  HDOA21M20D1 U1878 ( .A1(n2484), .A2(n1784), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n136), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n128) );
  HDAND2D1 U1879 ( .A1(n1805), .A2(n1734), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n935) );
  HDNAN2D1 U1880 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[10]), .Z(
        n1588) );
  HDOAI211D1 U1881 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[10]), .B(
        byp_alu_rs1_data_e[10]), .C(n1588), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n892) );
  HDNAN2D1 U1882 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[11]), .Z(
        n1589) );
  HDOAI211D1 U1883 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[11]), .B(
        byp_alu_rs1_data_e[11]), .C(n1589), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n881) );
  HDOAI22D1 U1884 ( .A1(n3383), .A2(n3096), .B1(n3165), .B2(n3498), .Z(n1590)
         );
  HDOAI22D1 U1885 ( .A1(n3264), .A2(n2456), .B1(n3184), .B2(n2704), .Z(n1591)
         );
  HDNOR2D1 U1886 ( .A1(n1590), .A2(n1591), .Z(n3104) );
  HDNAN2D1 U1887 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[25]), .Z(
        n1592) );
  HDOAI211D1 U1888 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[25]), .B(
        byp_alu_rs1_data_e[25]), .C(n1592), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n708) );
  HDOAI22D1 U1889 ( .A1(n3203), .A2(n2710), .B1(n3287), .B2(n2709), .Z(n1593)
         );
  HDOAI22D1 U1890 ( .A1(n3358), .A2(n2456), .B1(n3202), .B2(n2704), .Z(n1594)
         );
  HDNOR2D1 U1891 ( .A1(n1593), .A2(n1594), .Z(n3269) );
  HDNAN2D1 U1892 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[41]), .Z(
        n1595) );
  HDOAI211D1 U1893 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[41]), .B(
        byp_alu_rs1_data_e[41]), .C(n1595), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n408) );
  HDNOR2M1D1 U1894 ( .A1(byp_alu_rs1_data_e[12]), .A2(ecl_shft_enshift_e_l), 
        .Z(n3529) );
  HDNOR2M1D1 U1895 ( .A1(byp_alu_rs1_data_e[7]), .A2(ecl_shft_enshift_e_l), 
        .Z(n3483) );
  HDOA21D1 U1896 ( .A1(n2275), .A2(n2177), .B(n1871), .Z(n2459) );
  HDNOR2M1D1 U1897 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n662), 
        .A2(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n651), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n649) );
  HDOA22DL U1898 ( .A1(n2696), .A2(n3567), .B1(n3566), .B2(n3565), .Z(n1596)
         );
  HDNAN2D1 U1899 ( .A1(n2662), .A2(byp_alu_rs1_data_e[63]), .Z(n1597) );
  HDOAI211D1 U1900 ( .A1(n1744), .A2(n3568), .B(n1596), .C(n1597), .Z(n2264)
         );
  HDNAN2D1 U1901 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[5]), .Z(n1598) );
  HDOAI211D1 U1902 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[5]), .B(
        byp_alu_rs1_data_e[5]), .C(n1598), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n938) );
  HDOA21M20D1 U1903 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n886), 
        .A2(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n999), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n881), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n873) );
  HDAOI22D1 U1904 ( .A1(n3010), .A2(ecl_shft_shift4_e[3]), .B1(
        ecl_shft_shift4_e[1]), .B2(n3084), .Z(n1599) );
  HDNAN2D1 U1905 ( .A1(n3011), .A2(ecl_shft_shift4_e[0]), .Z(n1600) );
  HDOA211D1 U1906 ( .A1(n3119), .A2(n2707), .B(n1599), .C(n1600), .Z(n3057) );
  HDAOI21M10D1 U1907 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n764), 
        .A2(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n839), .B(n2315), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n761) );
  HDNAN2M1D1 U1908 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n725), 
        .A2(n2134), .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n604) );
  HDNAN2D1 U1909 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[26]), .Z(
        n1601) );
  HDOAI211D1 U1910 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[26]), .B(
        byp_alu_rs1_data_e[26]), .C(n1601), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n695) );
  HDOAI22D1 U1911 ( .A1(n3203), .A2(n2705), .B1(n3394), .B2(n3165), .Z(n1602)
         );
  HDOAI22D1 U1912 ( .A1(n3287), .A2(n2704), .B1(n3202), .B2(n2456), .Z(n1603)
         );
  HDNOR2D1 U1913 ( .A1(n1602), .A2(n1603), .Z(n3185) );
  HDNAN2D1 U1914 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[28]), .Z(
        n1604) );
  HDOAI211D1 U1915 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[28]), .B(
        byp_alu_rs1_data_e[28]), .C(n1604), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n669) );
  HDOAI22D1 U1916 ( .A1(n2205), .A2(n2456), .B1(n3332), .B2(n2704), .Z(n1605)
         );
  HDOAI22D1 U1917 ( .A1(n3224), .A2(n2710), .B1(n3223), .B2(n2709), .Z(n1606)
         );
  HDNOR2D1 U1918 ( .A1(n1605), .A2(n1606), .Z(n3291) );
  HDNAN2D1 U1919 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[33]), .Z(
        n1607) );
  HDOAI211D1 U1920 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[33]), .B(
        byp_alu_rs1_data_e[33]), .C(n1607), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n544) );
  HDNOR2M1D1 U1921 ( .A1(byp_alu_rs1_data_e[43]), .A2(n2588), .Z(n2125) );
  HDEXOR2DL U1922 ( .A1(byp_alu_rs1_data_e[63]), .A2(alu_addsub_rs2_data[63]), 
        .Z(n2266) );
  HDNAN2D1 U1923 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n977), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n1010), .Z(n1608) );
  HDEXNOR2DL U1924 ( .A1(alu_addsub_rs2_data[0]), .A2(n1608), .Z(
        alu_adder_out[0]) );
  HDEXOR2DL U1925 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[2]), .Z(
        n1609) );
  HDINVDL U1926 ( .A(n1772), .Z(n1610) );
  HDNAN2D1 U1927 ( .A1(n1609), .A2(n1767), .Z(n1611) );
  HDOAI211D1 U1928 ( .A1(n1609), .A2(n1610), .B(n1769), .C(n1611), .Z(n2780)
         );
  HDNAN2D1 U1929 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n1006), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n951), .Z(n1612) );
  HDAOI21D1 U1930 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n953), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n961), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n954), .Z(n1613) );
  HDEXOR2DL U1931 ( .A1(n1612), .A2(n1613), .Z(alu_adder_out[4]) );
  HDAOI22M10D1 U1932 ( .B1(n2695), .B2(n3120), .A1(n3566), .A2(n1756), .Z(
        n1614) );
  HDOAI211D1 U1933 ( .A1(n2685), .A2(n3498), .B(n3347), .C(n1614), .Z(n2818)
         );
  HDNAN2D1 U1934 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[17]), .Z(
        n1615) );
  HDOAI211D1 U1935 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[17]), .B(
        byp_alu_rs1_data_e[17]), .C(n1615), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n804) );
  HDNOR2M1D1 U1936 ( .A1(byp_alu_rs1_data_e[42]), .A2(n2396), .Z(n2194) );
  HDAO21D1 U1937 ( .A1(ecl_shft_shift4_e[0]), .A2(n3528), .B(n3527), .Z(n3548)
         );
  HDNAN2D1 U1938 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[6]), .Z(n1616) );
  HDOAI211D1 U1939 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[6]), .B(
        byp_alu_rs1_data_e[6]), .C(n1616), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n933) );
  HDNAN2M1D1 U1940 ( .A1(n1999), .A2(n1772), .Z(n2540) );
  HDOA21M20D1 U1941 ( .A1(n2465), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n896), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n903), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n895) );
  HDOA21M20DL U1942 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n886), 
        .A2(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n863), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n866), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n862) );
  HDNAN2M1DL U1943 ( .A1(n1732), .A2(n1772), .Z(n2554) );
  HDAOI22D1 U1944 ( .A1(n2572), .A2(n1772), .B1(n1794), .B2(n1767), .Z(n1617)
         );
  HDNAN2D1 U1945 ( .A1(n1769), .A2(n1617), .Z(n2571) );
  HDNAN2M1D1 U1946 ( .A1(n2162), .A2(n1772), .Z(n2640) );
  HDAOI22D1 U1947 ( .A1(n2111), .A2(n1767), .B1(n1772), .B2(n2533), .Z(n1618)
         );
  HDNAN2D1 U1948 ( .A1(n1769), .A2(n1618), .Z(n1619) );
  HDAOI22D1 U1949 ( .A1(byp_alu_rs2_data_e[23]), .A2(n2683), .B1(
        byp_alu_rs1_data_e[23]), .B2(n1619), .Z(n2532) );
  HDNAN2M1D1 U1950 ( .A1(n2130), .A2(n1772), .Z(n2625) );
  HDAOI22M20D1 U1951 ( .B1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n649), 
        .B2(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n689), .A1(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n651), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n665), .Z(n1620) );
  HDOAI211D1 U1952 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n739), 
        .A2(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n647), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n652), .C(n1620), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n646) );
  HDOAI22D1 U1953 ( .A1(n3184), .A2(n2710), .B1(n3264), .B2(n2708), .Z(n1621)
         );
  HDOAI22D1 U1954 ( .A1(n3349), .A2(n2456), .B1(n3183), .B2(n2704), .Z(n1622)
         );
  HDNOR2D1 U1955 ( .A1(n1621), .A2(n1622), .Z(n3245) );
  HDINVDL U1956 ( .A(n1772), .Z(n1623) );
  HDNAN2D1 U1957 ( .A1(n2151), .A2(n1767), .Z(n1624) );
  HDOAI211D1 U1958 ( .A1(n2151), .A2(n1623), .B(n1769), .C(n1624), .Z(n2445)
         );
  HDNAN2M1D1 U1959 ( .A1(n2186), .A2(n1772), .Z(n2076) );
  HDNOR2M1D1 U1960 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n227), 
        .A2(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n195), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n193) );
  HDAOI22M10D1 U1961 ( .B1(ecl_shft_shift4_e[3]), .B2(n2126), .A1(n2456), .A2(
        n2264), .Z(n1625) );
  HDOAI21M20DL U1962 ( .A1(n1625), .A2(n2263), .B(ecl_shft_shift1_e[0]), .Z(
        n1626) );
  HDOAI21M20DL U1963 ( .A1(n3571), .A2(ecl_shft_shift1_e[1]), .B(n1626), .Z(
        n2258) );
  HDOAI21M10D1 U1964 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n1009), 
        .A2(n2475), .B(n1872), .Z(n1627) );
  HDNAN2M1D1 U1965 ( .A1(n1737), .A2(n1738), .Z(n1628) );
  HDEXNOR2DL U1966 ( .A1(n1628), .A2(n1627), .Z(alu_adder_out[2]) );
  HDNAN2D1 U1967 ( .A1(n1805), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n938), .Z(n1629) );
  HDAOI21DL U1968 ( .A1(n1734), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n961), .B(n2477), .Z(n1630)
         );
  HDEXOR2DL U1969 ( .A1(n1629), .A2(n1630), .Z(alu_adder_out[5]) );
  HDOAI222D1 U1970 ( .A1(n2894), .A2(n1783), .B1(n2882), .B2(n2686), .C1(n2924), .C2(n1789), .Z(n1631) );
  HDAOI21M10D1 U1971 ( .A1(n2904), .A2(n2692), .B(n1631), .Z(n2543) );
  HDNAN2D1 U1972 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n995), .A2(
        n2177), .Z(n1632) );
  HDEXNOR2DL U1973 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n839), 
        .A2(n1632), .Z(alu_adder_out[15]) );
  HDAOI22D1 U1974 ( .A1(n3099), .A2(ecl_shft_shift4_e[2]), .B1(
        ecl_shft_shift4_e[1]), .B2(n3043), .Z(n1633) );
  HDNAN2D1 U1975 ( .A1(ecl_shft_shift4_e[0]), .A2(n2981), .Z(n1634) );
  HDOA211D1 U1976 ( .A1(n3158), .A2(n2710), .B(n1633), .C(n1634), .Z(n3025) );
  HDOA21M10DL U1977 ( .A2(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n464), 
        .A1(n2431), .B(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n447), .Z(
        n2419) );
  HDNAN2M1D1 U1978 ( .A1(n2689), .A2(byp_alu_rs2_data_e[41]), .Z(n2085) );
  HDOAI222D1 U1979 ( .A1(n3368), .A2(n3533), .B1(n3377), .B2(n3576), .C1(n2359), .C2(n1789), .Z(n1635) );
  HDNOR2D1 U1980 ( .A1(n3387), .A2(n3563), .Z(n1636) );
  HDNOR3D1 U1981 ( .A1(n1636), .A2(n1635), .A3(n2055), .Z(n2050) );
  HDNAN2M1D1 U1982 ( .A1(n2125), .A2(n2490), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n25) );
  HDNAN2M1D1 U1983 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n361), 
        .A2(n2013), .Z(n2398) );
  HDNOR4D1 U1984 ( .A1(n1900), .A2(n1901), .A3(n1902), .A4(n1899), .Z(n1637)
         );
  HDNAN2D1 U1985 ( .A1(n1765), .A2(byp_alu_rs2_data_e[46]), .Z(n1638) );
  HDOAI21D1 U1986 ( .A1(n1637), .A2(ecl_alu_out_sel_shift_e_l), .B(n1638), .Z(
        n1898) );
  HDMUXB2DL U1987 ( .A0(n1772), .A1(n1767), .SL(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_23_), .Z(n1639) );
  HDOA21M20D1 U1988 ( .A1(n1769), .A2(n1639), .B(byp_alu_rs1_data_e[55]), .Z(
        n2029) );
  HDNAN3M1DL U1989 ( .A1(n2349), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n158), .A3(n1785), .Z(n2356) );
  HDOAI21DL U1990 ( .A1(n2703), .A2(byp_alu_rs1_data_e[60]), .B(n1769), .Z(
        n1640) );
  HDNAN2D1 U1991 ( .A1(n2645), .A2(n1772), .Z(n1641) );
  HDNAN3DL U1992 ( .A1(n1641), .A2(n2644), .A3(n1769), .Z(n1642) );
  HDAO22DL U1993 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_28_), 
        .A2(n1640), .B1(byp_alu_rs1_data_e[60]), .B2(n1642), .Z(n2650) );
  HDNAN2D1 U1994 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[16]), .Z(
        n1643) );
  HDOAI211D1 U1995 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[16]), .B(
        byp_alu_rs1_data_e[16]), .C(n1643), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n825) );
  HDOA21M20D1 U1996 ( .A1(n2473), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n985), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n708), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n700) );
  HDAOI211D1 U1997 ( .A1(byp_alu_rs1_data_e[43]), .A2(n2699), .B(n2574), .C(
        n3375), .Z(n1644) );
  HDNOR2D1 U1998 ( .A1(n2456), .A2(n1644), .Z(n2575) );
  HDNOR2M1D1 U1999 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n363), 
        .A2(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n331), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n329) );
  HDAO22DL U2000 ( .A1(n2203), .A2(byp_alu_rs1_data_e[60]), .B1(n3536), .B2(
        n3529), .Z(n2549) );
  HDNAN2M1D1 U2001 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n905), 
        .A2(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n896), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n894) );
  HDNAN2D1 U2002 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n886), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n852), .Z(n1645) );
  HDOA211DL U2003 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n854), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n866), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n855), .C(n1645), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n851) );
  HDOAI22D1 U2004 ( .A1(n3200), .A2(n2456), .B1(n3284), .B2(n2704), .Z(n1646)
         );
  HDOAI22D1 U2005 ( .A1(n3319), .A2(n2708), .B1(n3199), .B2(n2710), .Z(n1647)
         );
  HDNOR2D1 U2006 ( .A1(n1646), .A2(n1647), .Z(n3270) );
  HDEXOR2DL U2007 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[36]), .Z(
        n1648) );
  HDMUXB2DL U2008 ( .A0(n1772), .A1(n1767), .SL(n1648), .Z(n2247) );
  HDMUXB2DL U2009 ( .A0(n1772), .A1(n1767), .SL(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_15_), .Z(n1649) );
  HDAOI21D1 U2010 ( .A1(n1649), .A2(n1769), .B(n3568), .Z(n2387) );
  HDNAN2M1D1 U2011 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_19_), 
        .A2(n1772), .Z(n2092) );
  HDNAN2D1 U2012 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[52]), .Z(
        n1650) );
  HDOAI211D1 U2013 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[52]), .B(
        byp_alu_rs1_data_e[52]), .C(n1650), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n209) );
  HDNAN2D1 U2014 ( .A1(n2483), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n117), .Z(n1651) );
  HDOAI211D1 U2015 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n128), 
        .A2(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n97), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n102), .C(n1651), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n96) );
  HDNOR2D1 U2016 ( .A1(n3574), .A2(n2702), .Z(n1652) );
  HDNOR2D1 U2017 ( .A1(n3575), .A2(n3576), .Z(n1653) );
  HDNOR3D1 U2018 ( .A1(n1653), .A2(n3577), .A3(n1652), .Z(n2262) );
  HDNAN2D1 U2019 ( .A1(n1872), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n1009), .Z(n1654) );
  HDEXOR2DL U2020 ( .A1(n1654), .A2(n2475), .Z(alu_adder_out[1]) );
  HDOAI22D1 U2021 ( .A1(n3560), .A2(n2802), .B1(n2774), .B2(n2702), .Z(n1655)
         );
  HDOAI22D1 U2022 ( .A1(n1783), .A2(n2792), .B1(n2817), .B2(n3561), .Z(n1656)
         );
  HDNOR3D1 U2023 ( .A1(n2779), .A2(n1655), .A3(n1656), .Z(n2784) );
  HDEXOR2DL U2024 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[3]), .Z(
        n1657) );
  HDINVDL U2025 ( .A(n1772), .Z(n1658) );
  HDNAN2D1 U2026 ( .A1(n1657), .A2(n1767), .Z(n1659) );
  HDOAI211D1 U2027 ( .A1(n1657), .A2(n1658), .B(n1769), .C(n1659), .Z(n2797)
         );
  HDINVDL U2028 ( .A(n1772), .Z(n1660) );
  HDNAN2D1 U2029 ( .A1(n2000), .A2(n1767), .Z(n1661) );
  HDOAI211D1 U2030 ( .A1(n2000), .A2(n1660), .B(n1769), .C(n1661), .Z(n2812)
         );
  HDAOI21D1 U2031 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n935), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n961), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n936), .Z(n1662) );
  HDNAN2M1D1 U2032 ( .A1(n2108), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n933), .Z(n1663) );
  HDEXOR2DL U2033 ( .A1(n1663), .A2(n1662), .Z(alu_adder_out[6]) );
  HDOAI21D1 U2034 ( .A1(n2703), .A2(byp_alu_rs1_data_e[9]), .B(n1769), .Z(
        n1664) );
  HDNAN3D1 U2035 ( .A1(n1769), .A2(n2541), .A3(n2540), .Z(n1665) );
  HDAO222D1 U2036 ( .A1(n1664), .A2(n1998), .B1(n1665), .B2(
        byp_alu_rs1_data_e[9]), .C1(n2683), .C2(byp_alu_rs2_data_e[9]), .Z(
        n2539) );
  HDINVDL U2037 ( .A(n1772), .Z(n1666) );
  HDNAN2D1 U2038 ( .A1(n2274), .A2(n1767), .Z(n1667) );
  HDOAI211D1 U2039 ( .A1(n2274), .A2(n1666), .B(n1769), .C(n1667), .Z(n2899)
         );
  HDOAI21D1 U2040 ( .A1(n2703), .A2(byp_alu_rs1_data_e[16]), .B(n1769), .Z(
        n1668) );
  HDNAN3D1 U2041 ( .A1(n1769), .A2(n2555), .A3(n2554), .Z(n1669) );
  HDAO222D1 U2042 ( .A1(n1668), .A2(n1731), .B1(n1669), .B2(
        byp_alu_rs1_data_e[16]), .C1(n2683), .C2(byp_alu_rs2_data_e[16]), .Z(
        n2553) );
  HDNAN2D1 U2043 ( .A1(n1793), .A2(n1815), .Z(n1670) );
  HDNAN2D1 U2044 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n813), .A2(
        n1670), .Z(n1671) );
  HDOAI211D1 U2045 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n813), 
        .A2(n1670), .B(n1785), .C(n1671), .Z(n2564) );
  HDEXOR2DL U2046 ( .A1(byp_alu_rs2_data_e[19]), .A2(ifu_exu_invert_d), .Z(
        n1672) );
  HDINVDL U2047 ( .A(n1772), .Z(n1673) );
  HDNAN2D1 U2048 ( .A1(n1672), .A2(n1767), .Z(n1674) );
  HDOAI211D1 U2049 ( .A1(n1672), .A2(n1673), .B(n1769), .C(n1674), .Z(n3052)
         );
  HDOAI21D1 U2050 ( .A1(n2703), .A2(byp_alu_rs1_data_e[21]), .B(n1769), .Z(
        n1675) );
  HDNAN3D1 U2051 ( .A1(n1769), .A2(n2641), .A3(n2640), .Z(n1676) );
  HDAO222D1 U2052 ( .A1(n1675), .A2(n2162), .B1(n1676), .B2(
        byp_alu_rs1_data_e[21]), .C1(n2683), .C2(byp_alu_rs2_data_e[21]), .Z(
        n2639) );
  HDOAI21D1 U2053 ( .A1(n2703), .A2(byp_alu_rs1_data_e[24]), .B(n1769), .Z(
        n1677) );
  HDNAN3D1 U2054 ( .A1(n1769), .A2(n2626), .A3(n2625), .Z(n1678) );
  HDAO222D1 U2055 ( .A1(n1677), .A2(n2130), .B1(n1678), .B2(
        byp_alu_rs1_data_e[24]), .C1(n2683), .C2(byp_alu_rs2_data_e[24]), .Z(
        n2624) );
  HDOAI22D1 U2056 ( .A1(n3246), .A2(n3561), .B1(n1789), .B2(n3245), .Z(n3189)
         );
  HDOA22DL U2057 ( .A1(n3560), .A2(n3300), .B1(n3299), .B2(n3563), .Z(n1679)
         );
  HDOA22DL U2058 ( .A1(n3292), .A2(n2702), .B1(n3291), .B2(n3533), .Z(n1680)
         );
  HDNAN4D1 U2059 ( .A1(n2437), .A2(n2439), .A3(n1679), .A4(n1680), .Z(n2438)
         );
  HDNAN2M1D1 U2060 ( .A1(n2689), .A2(byp_alu_rs2_data_e[35]), .Z(n1947) );
  HDOAI21D1 U2061 ( .A1(n2703), .A2(byp_alu_rs1_data_e[37]), .B(n1769), .Z(
        n1681) );
  HDINVDL U2062 ( .A(n1772), .Z(n1682) );
  HDNAN2D1 U2063 ( .A1(n1934), .A2(n1767), .Z(n1683) );
  HDOAI211D1 U2064 ( .A1(n1934), .A2(n1682), .B(n1769), .C(n1683), .Z(n1684)
         );
  HDAO22DL U2065 ( .A1(n1967), .A2(n1681), .B1(byp_alu_rs1_data_e[37]), .B2(
        n1684), .Z(n1929) );
  HDNOR2M1D1 U2066 ( .A1(n1785), .A2(n2430), .Z(n1753) );
  HDOAI21D1 U2067 ( .A1(byp_alu_rs1_data_e[40]), .A2(n2703), .B(n1769), .Z(
        n1685) );
  HDNAN2D1 U2068 ( .A1(n1685), .A2(n2120), .Z(n1686) );
  HDEXOR2DL U2069 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[40]), .Z(
        n1687) );
  HDMUXB2DL U2070 ( .A0(n1772), .A1(n1767), .SL(n1687), .Z(n1688) );
  HDAOI32D1 U2071 ( .A1(n1769), .A2(n1686), .A3(n1688), .B1(n3346), .B2(n1686), 
        .Z(n2499) );
  HDOAI21D1 U2072 ( .A1(byp_alu_rs1_data_e[41]), .A2(n2703), .B(n1769), .Z(
        n1689) );
  HDAOI31D1 U2073 ( .A1(n2077), .A2(n1769), .A3(n2076), .B(n3355), .Z(n1690)
         );
  HDAOI21D1 U2074 ( .A1(n2186), .A2(n1689), .B(n1690), .Z(n2087) );
  HDNAN3D1 U2075 ( .A1(n1769), .A2(n2054), .A3(n2053), .Z(n1691) );
  HDEXOR2DL U2076 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[42]), .Z(
        n1692) );
  HDOAI21D1 U2077 ( .A1(n2703), .A2(byp_alu_rs1_data_e[42]), .B(n1769), .Z(
        n1693) );
  HDAOI22D1 U2078 ( .A1(byp_alu_rs1_data_e[42]), .A2(n1691), .B1(n1692), .B2(
        n1693), .Z(n2051) );
  HDNAN3D1 U2079 ( .A1(n1769), .A2(n2044), .A3(n2043), .Z(n1694) );
  HDEXOR2DL U2080 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[43]), .Z(
        n1695) );
  HDOAI21D1 U2081 ( .A1(n2703), .A2(byp_alu_rs1_data_e[43]), .B(n1769), .Z(
        n1696) );
  HDAOI22D1 U2082 ( .A1(byp_alu_rs1_data_e[43]), .A2(n1694), .B1(n1695), .B2(
        n1696), .Z(n2041) );
  HDOAI21D1 U2083 ( .A1(n2703), .A2(byp_alu_rs1_data_e[45]), .B(n1769), .Z(
        n1697) );
  HDOAI21M20DL U2084 ( .A1(n1769), .A2(n1912), .B(byp_alu_rs1_data_e[45]), .Z(
        n1698) );
  HDOAI21M20DL U2085 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_13_), 
        .A2(n1697), .B(n1698), .Z(n1913) );
  HDOAI21D1 U2086 ( .A1(n2703), .A2(byp_alu_rs1_data_e[46]), .B(n1769), .Z(
        n1699) );
  HDINVDL U2087 ( .A(n1772), .Z(n1700) );
  HDNAN2D1 U2088 ( .A1(n1904), .A2(n1767), .Z(n1701) );
  HDOAI211D1 U2089 ( .A1(n1904), .A2(n1700), .B(n1769), .C(n1701), .Z(n1702)
         );
  HDAO22DL U2090 ( .A1(n2104), .A2(n1699), .B1(byp_alu_rs1_data_e[46]), .B2(
        n1702), .Z(n1903) );
  HDNOR2M1D1 U2091 ( .A1(n1785), .A2(n2392), .Z(n1739) );
  HDOAI21D1 U2092 ( .A1(byp_alu_rs1_data_e[48]), .A2(n2703), .B(n1769), .Z(
        n1703) );
  HDNAN2D1 U2093 ( .A1(n1703), .A2(n1977), .Z(n1704) );
  HDEXOR2DL U2094 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[48]), .Z(
        n1705) );
  HDMUXB2DL U2095 ( .A0(n1772), .A1(n1767), .SL(n1705), .Z(n1706) );
  HDAOI32D1 U2096 ( .A1(n1769), .A2(n1704), .A3(n1706), .B1(n3414), .B2(n1704), 
        .Z(n2667) );
  HDNOR2M1D1 U2097 ( .A1(byp_alu_rs2_data_e[51]), .A2(n2689), .Z(n2100) );
  HDOAI21D1 U2098 ( .A1(n2703), .A2(byp_alu_rs1_data_e[53]), .B(n1769), .Z(
        n1707) );
  HDOAI21M20DL U2099 ( .A1(n1769), .A2(n1917), .B(byp_alu_rs1_data_e[53]), .Z(
        n1708) );
  HDOAI21M20DL U2100 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_21_), 
        .A2(n1707), .B(n1708), .Z(n1922) );
  HDNAN4M1D1 U2101 ( .A1(n2313), .A2(n1785), .A3(n2312), .A4(n2311), .Z(n2024)
         );
  HDNOR2D1 U2102 ( .A1(n3519), .A2(n3561), .Z(n1709) );
  HDNOR3D1 U2103 ( .A1(n1709), .A2(n2354), .A3(n2353), .Z(n1710) );
  HDOAI21D1 U2104 ( .A1(n2591), .A2(n3533), .B(n1710), .Z(n2350) );
  HDOAI21D1 U2105 ( .A1(n2703), .A2(byp_alu_rs1_data_e[57]), .B(n1769), .Z(
        n1711) );
  HDINVDL U2106 ( .A(n1772), .Z(n1712) );
  HDNAN2D1 U2107 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_25_), 
        .A2(n1767), .Z(n1713) );
  HDOAI211D1 U2108 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_25_), 
        .A2(n1712), .B(n1769), .C(n1713), .Z(n1714) );
  HDAO22DL U2109 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_25_), 
        .A2(n1711), .B1(byp_alu_rs1_data_e[57]), .B2(n1714), .Z(n2374) );
  HDOAI22D1 U2110 ( .A1(n3508), .A2(n3533), .B1(n3534), .B2(n1789), .Z(n1715)
         );
  HDNOR2D1 U2111 ( .A1(n3518), .A2(n1783), .Z(n1716) );
  HDNOR3D1 U2112 ( .A1(n1716), .A2(n1715), .A3(n2601), .Z(n2593) );
  HDNOR2M1D1 U2113 ( .A1(byp_alu_rs2_data_e[60]), .A2(n2689), .Z(n2652) );
  HDOAI21D1 U2114 ( .A1(n2703), .A2(byp_alu_rs1_data_e[63]), .B(n1769), .Z(
        n1717) );
  HDOAI211D1 U2115 ( .A1(alu_addsub_rs2_data[63]), .A2(n2703), .B(n1769), .C(
        n2257), .Z(n1718) );
  HDAO222D1 U2116 ( .A1(n1717), .A2(alu_addsub_rs2_data[63]), .B1(n1718), .B2(
        byp_alu_rs1_data_e[63]), .C1(n3579), .C2(byp_alu_rs2_data_e[63]), .Z(
        n2256) );
  HDNOR3D1 U2117 ( .A1(n2535), .A2(n2534), .A3(n2536), .Z(n1719) );
  HDNAN2M1D1 U2118 ( .A1(ecl_alu_out_sel_shift_e_l), .A2(n2530), .Z(n1720) );
  HDOAI211D1 U2119 ( .A1(ecl_alu_out_sel_shift_e_l), .A2(n1719), .B(n2529), 
        .C(n1720), .Z(alu_byp_rd_data_e[23]) );
  HDNOR2D1 U2120 ( .A1(n2399), .A2(n2400), .Z(n1721) );
  HDNAN4D1 U2121 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n362), .A2(
        n1785), .A3(n2412), .A4(n2398), .Z(n1722) );
  HDOAI211D1 U2122 ( .A1(n2397), .A2(n2398), .B(n1721), .C(n1722), .Z(
        alu_byp_rd_data_e[44]) );
  HDOAI22M10D1 U2123 ( .A1(n3562), .A2(n3204), .B1(n3205), .B2(n3576), .Z(
        n3187) );
  HDOA22D2 U2124 ( .A1(n3294), .A2(n2702), .B1(n3293), .B2(n3533), .Z(n1954)
         );
  HDINVDL U2125 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n532), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n530) );
  HDAOI211D4 U2126 ( .A1(ecl_shft_shift4_e[3]), .A2(n3467), .B(n2618), .C(
        n2619), .Z(n2591) );
  HDINVD2 U2127 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n840), .Z(
        n1723) );
  HDINVBD2 U2128 ( .A(n1723), .Z(n1724) );
  HDNAN2D8 U2129 ( .A1(n2454), .A2(byp_alu_rs2_data_e[4]), .Z(n1773) );
  HDOAI22M10D1 U2130 ( .A1(n3579), .A2(n1725), .B1(n2243), .B2(
        ecl_alu_out_sel_shift_e_l), .Z(n2242) );
  HDINVDL U2131 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n798), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n992) );
  HDOA211D1 U2132 ( .A1(n1726), .A2(n1727), .B(n1728), .C(n1729), .Z(n2773) );
  HDOA22D1 U2133 ( .A1(n2802), .A2(n3561), .B1(n2774), .B2(n3576), .Z(n1728)
         );
  HDOA222D4 U2134 ( .A1(n3563), .A2(n2792), .B1(n2702), .B2(n2766), .C1(n3560), 
        .C2(n2785), .Z(n1729) );
  HDNAN2D1 U2135 ( .A1(n2105), .A2(byp_alu_rs1_data_e[30]), .Z(n1730) );
  HDNAN2D1 U2136 ( .A1(n2105), .A2(byp_alu_rs1_data_e[30]), .Z(n3402) );
  HDAND2D2 U2137 ( .A1(n3460), .A2(n3459), .Z(n3531) );
  HDEXOR2D1 U2138 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[16]), .Z(
        n1732) );
  HDEXOR2DL U2139 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[16]), .Z(
        n1731) );
  HDBUFD1 U2140 ( .A(n2785), .Z(n1733) );
  HDINVDL U2141 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n752), .Z(
        n2316) );
  HDNOR2DL U2142 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n950), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n959), .Z(n1734) );
  HDNOR2D1 U2143 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n950), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n959), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n944) );
  HDNAN2D1 U2144 ( .A1(n2756), .A2(ecl_alu_log_sel_xor_e), .Z(n1735) );
  HDINVBD16 U2145 ( .A(n1735), .Z(n1772) );
  HDNAN2DL U2146 ( .A1(n2357), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n778), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n608) );
  HDOAI211D2 U2147 ( .A1(n2788), .A2(n1773), .B(n2961), .C(n2787), .Z(n2981)
         );
  HDAND3D1 U2148 ( .A1(n1798), .A2(n1799), .A3(n1796), .Z(n1736) );
  HDAND3D1 U2149 ( .A1(n1798), .A2(n1799), .A3(n1796), .Z(n1737) );
  HDOR2D1 U2150 ( .A1(n1732), .A2(byp_alu_rs1_data_e[16]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n994) );
  HDBUFDL U2151 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n966), .Z(
        n1738) );
  HDNAN3D1 U2152 ( .A1(n2376), .A2(n2384), .A3(n1739), .Z(n2378) );
  HDNAN2M1D2 U2153 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n191), 
        .A2(n2190), .Z(n2218) );
  HDAO21D2 U2154 ( .A1(n2470), .A2(n3282), .B(n1740), .Z(n3417) );
  HDNOR2D1 U2155 ( .A1(n2527), .A2(n2528), .Z(n2526) );
  HDNAN3D2 U2156 ( .A1(n2415), .A2(n2419), .A3(n1753), .Z(n2416) );
  HDINVD12 U2157 ( .A(byp_alu_rs2_data_e[5]), .Z(n1741) );
  HDINVD4 U2158 ( .A(n1741), .Z(n1742) );
  HDOR2D4 U2159 ( .A1(n2506), .A2(ecl_shft_enshift_e_l), .Z(n1743) );
  HDOR2D4 U2160 ( .A1(n2506), .A2(ecl_shft_enshift_e_l), .Z(n1744) );
  HDOAI22M10D1 U2161 ( .A1(n1745), .A2(n1779), .B1(n3406), .B2(n3576), .Z(
        n1900) );
  HDNAN2D6 U2162 ( .A1(n2454), .A2(byp_alu_rs2_data_e[4]), .Z(n2675) );
  HDNAN2DL U2163 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n990), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n773), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n607) );
  HDOAI22D2 U2164 ( .A1(n2300), .A2(n2709), .B1(n2205), .B2(n2710), .Z(n2364)
         );
  HDOA21D1 U2165 ( .A1(n1743), .A2(n3448), .B(n3447), .Z(n2107) );
  HDOA21M20D2 U2166 ( .A1(n2088), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n397), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n404), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n396) );
  HDOAI21M10D1 U2167 ( .A1(byp_alu_rs1_data_e[41]), .A2(ecl_shft_op32_e), .B(
        n2678), .Z(n3139) );
  HDINVD1 U2168 ( .A(byp_alu_rs1_data_e[41]), .Z(n3355) );
  HDNOR2M1D2 U2169 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n994), 
        .A2(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n837), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n814) );
  HDINVD12 U2170 ( .A(n2695), .Z(n2693) );
  HDOR2D2 U2171 ( .A1(n3525), .A2(n1783), .Z(n1835) );
  HDINVBD4 U2172 ( .A(ifu_exu_invert_d), .Z(n1800) );
  HDINVBD4 U2173 ( .A(ifu_exu_invert_d), .Z(n1971) );
  HDINVBD2 U2174 ( .A(ifu_exu_invert_d), .Z(n1970) );
  HDINVD2 U2175 ( .A(ifu_exu_invert_d), .Z(n1873) );
  HDNOR2D2 U2176 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I2_20_), 
        .A2(byp_alu_rs1_data_e[20]), .Z(n1748) );
  HDOAI22DL U2177 ( .A1(n3296), .A2(n2710), .B1(n3220), .B2(n2707), .Z(n3091)
         );
  HDOAI22DL U2178 ( .A1(n3284), .A2(n2710), .B1(n3200), .B2(n2707), .Z(n3083)
         );
  HDINVD8 U2179 ( .A(n2684), .Z(n2685) );
  HDOA21M20D2 U2180 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n3), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n227), .B(n2467), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n226) );
  HDNAN2D2 U2181 ( .A1(n2653), .A2(byp_alu_rs1_data_e[20]), .Z(n3315) );
  HDNAN2D1 U2182 ( .A1(n2653), .A2(byp_alu_rs1_data_e[24]), .Z(n3347) );
  HDINVD4 U2183 ( .A(n2693), .Z(n2697) );
  HDINVD4 U2184 ( .A(n2696), .Z(n1786) );
  HDINVD16 U2185 ( .A(n2679), .Z(n2676) );
  HDOAI21M20DL U2186 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n793), 
        .A2(n2357), .B(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n778), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n776) );
  HDNAN2DL U2187 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n792), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n766), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n764) );
  HDNAN3D2 U2188 ( .A1(n2607), .A2(n2606), .A3(n2608), .Z(
        alu_byp_rd_data_e[62]) );
  HDEXOR2DL U2189 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[21]), .Z(
        n2162) );
  HDOAI22M10D1 U2190 ( .A1(ecl_shft_shift4_e[2]), .A2(n3539), .B1(n1749), .B2(
        n2589), .Z(n3506) );
  HDOAI22M10D1 U2191 ( .A1(n1751), .A2(n1986), .B1(n1750), .B2(n3524), .Z(
        n2209) );
  HDOA22D2 U2192 ( .A1(n1789), .A2(n2792), .B1(n2755), .B2(n3578), .Z(n2671)
         );
  HDAO21M20D1 U2193 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n90), 
        .A2(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n55), .B(n1752), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n54) );
  HDNAN2D2 U2194 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n432), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n363), .Z(n2375) );
  HDOA211D1 U2195 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n472), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n437), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n442), .C(n2337), .Z(n2338)
         );
  HDNAN2DL U2196 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n306), .A2(
        n2489), .Z(n2392) );
  HDAOI211D4 U2197 ( .A1(n3139), .A2(n1782), .B(n3176), .C(n3138), .Z(n3328)
         );
  HDEXOR2D1 U2198 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[32]), .Z(
        alu_addsub_rs2_data[32]) );
  HDINVD2 U2199 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n294), .Z(
        n1754) );
  HDINVD2 U2200 ( .A(n2478), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n294) );
  HDINVD1 U2201 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n816), .Z(
        n1755) );
  HDINVD2 U2202 ( .A(n2200), .Z(n2118) );
  HDINVD2 U2203 ( .A(n2118), .Z(n2109) );
  HDOR2D2 U2204 ( .A1(n2187), .A2(byp_alu_rs1_data_e[41]), .Z(n2486) );
  HDNAN2D2 U2205 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n587), .A2(
        n2486), .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n403) );
  HDINVDL U2206 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n432), .Z(
        n2089) );
  HDINVDL U2207 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n814), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n816) );
  HDOA22D4 U2208 ( .A1(n3343), .A2(n3561), .B1(n3342), .B2(n1789), .Z(n1930)
         );
  HDAOI21M10D1 U2209 ( .A1(n2011), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n342), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n343), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n341) );
  HDINVD32 U2210 ( .A(byp_alu_rs2_data_e[5]), .Z(n2158) );
  HDINVD12 U2211 ( .A(n3566), .Z(n3536) );
  HDOA22M20D1 U2212 ( .A1(byp_alu_rs2_data_e[32]), .A2(n1758), .B1(n1759), 
        .B2(n1757), .Z(n3279) );
  HDBUFD4 U2213 ( .A(n3417), .Z(n2657) );
  HDOAI21M20D2 U2214 ( .A1(byp_alu_rs1_data_e[59]), .A2(n2745), .B(n2676), .Z(
        n1760) );
  HDOR2D2 U2215 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_13_), .A2(
        byp_alu_rs1_data_e[45]), .Z(n2493) );
  HDEXOR2DL U2216 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[35]), .Z(
        n1945) );
  HDNOR3D2 U2217 ( .A1(n1910), .A2(n1908), .A3(n1911), .Z(n1761) );
  HDNOR2D1 U2218 ( .A1(n1909), .A2(n1762), .Z(n1907) );
  HDINVD2 U2219 ( .A(n1761), .Z(n1762) );
  HDOAI22D2 U2220 ( .A1(n3406), .A2(n3560), .B1(n1779), .B2(n3563), .Z(n1909)
         );
  HDINVD2 U2221 ( .A(n2121), .Z(n2122) );
  HDOA21M20D2 U2222 ( .A1(n2336), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n435), .B(n2338), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n430) );
  HDBUFD2 U2223 ( .A(n2506), .Z(n2200) );
  HDAOI211D2 U2224 ( .A1(ecl_shft_shift4_e[2]), .A2(n3520), .B(n3456), .C(
        n3444), .Z(n3471) );
  HDINVD1 U2225 ( .A(n1764), .Z(n1763) );
  HDOAI22M10D1 U2226 ( .A1(byp_alu_rs2_data_e[45]), .A2(n1763), .B1(n1907), 
        .B2(ecl_alu_out_sel_shift_e_l), .Z(n1906) );
  HDBUFD8 U2227 ( .A(n3417), .Z(n2658) );
  HDINVD20 U2228 ( .A(byp_alu_rs2_data_e[5]), .Z(n2360) );
  HDNOR2D1 U2229 ( .A1(n3578), .A2(n1795), .Z(n1766) );
  HDINVBD16 U2230 ( .A(n1766), .Z(n3561) );
  HDINVD2 U2231 ( .A(ecl_shft_shift1_e[3]), .Z(n1795) );
  HDOA211D2 U2232 ( .A1(n3431), .A2(n3566), .B(n1824), .C(n1825), .Z(n3539) );
  HDAND2D1 U2233 ( .A1(ecl_shft_lshift_e_l), .A2(ecl_shft_shift1_e[0]), .Z(
        n2503) );
  HDOR2D4 U2234 ( .A1(n2199), .A2(n2198), .Z(n1768) );
  HDNOR2D6 U2235 ( .A1(n2757), .A2(ecl_alu_out_sel_logic_e_l), .Z(n1767) );
  HDINVD1 U2236 ( .A(n3563), .Z(n1788) );
  HDNAN2D4 U2237 ( .A1(n3578), .A2(ecl_shft_shift1_e[1]), .Z(n3563) );
  HDINVD1 U2238 ( .A(n3533), .Z(n2687) );
  HDINVBD4 U2239 ( .A(n3546), .Z(n3533) );
  HDINVD1 U2240 ( .A(n3560), .Z(n2692) );
  HDNAN2D4 U2241 ( .A1(ecl_shft_lshift_e_l), .A2(ecl_shft_shift1_e[2]), .Z(
        n3560) );
  HDINVD8 U2242 ( .A(ecl_shft_shift4_e[3]), .Z(n2710) );
  HDNAN2D8 U2243 ( .A1(n2756), .A2(ecl_alu_log_sel_or_e), .Z(n1769) );
  HDNAN2D1 U2244 ( .A1(n1968), .A2(byp_alu_rs1_data_e[29]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n652) );
  HDINVBD4 U2245 ( .A(ecl_alu_out_sel_sum_e_l), .Z(n1785) );
  HDAND2D1 U2246 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n499), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n465), .Z(n1771) );
  HDINVD2 U2247 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n736), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n738) );
  HDINVD2 U2248 ( .A(ecl_shft_shift4_e[2]), .Z(n2708) );
  HDINVD2 U2249 ( .A(ecl_shft_shift4_e[2]), .Z(n2706) );
  HDINVD2 U2250 ( .A(ecl_shft_shift4_e[2]), .Z(n2709) );
  HDINVD2 U2251 ( .A(ecl_shft_shift4_e[2]), .Z(n2707) );
  HDEXOR2DL U2252 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[17]), .Z(
        n1794) );
  HDINVBD4 U2253 ( .A(n2503), .Z(n2702) );
  HDEXOR2DL U2254 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[0]), .Z(
        alu_addsub_rs2_data[0]) );
  HDEXNOR2DL U2255 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[0]), .Z(
        n2135) );
  HDINVD1 U2256 ( .A(n2466), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n498) );
  HDINVD1 U2257 ( .A(n1869), .Z(n1790) );
  HDOR2D1 U2258 ( .A1(alu_addsub_rs2_data[42]), .A2(byp_alu_rs1_data_e[42]), 
        .Z(n1869) );
  HDOR2D1 U2259 ( .A1(n3493), .A2(n2710), .Z(n1774) );
  HDINVD1 U2260 ( .A(n2491), .Z(n2192) );
  HDINVD1 U2261 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n344), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n583) );
  HDINVD8 U2262 ( .A(ecl_shft_shift4_e[1]), .Z(n2704) );
  HDINVBD4 U2263 ( .A(n3562), .Z(n1783) );
  HDAND2D1 U2264 ( .A1(n3578), .A2(ecl_shft_shift1_e[2]), .Z(n3562) );
  HDOR2D1 U2265 ( .A1(n2035), .A2(n2034), .Z(n1775) );
  HDOR2D4 U2266 ( .A1(n2207), .A2(byp_alu_rs2_data_e[4]), .Z(n1776) );
  HDOR2D1 U2267 ( .A1(n2246), .A2(n2245), .Z(n1777) );
  HDINVD8 U2268 ( .A(ecl_shft_shift4_e[0]), .Z(n2456) );
  HDOR2D4 U2269 ( .A1(n2506), .A2(ecl_shft_enshift_e_l), .Z(n1778) );
  HDINVBD2 U2270 ( .A(n3579), .Z(n2689) );
  HDNOR2D2 U2271 ( .A1(n3278), .A2(ecl_alu_sethi_inst_e), .Z(n3579) );
  HDOA21D1 U2272 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n694), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n708), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n695), .Z(n1780) );
  HDINVD12 U2273 ( .A(ecl_shft_op32_e), .Z(n2745) );
  HDNOR2D2 U2274 ( .A1(n1878), .A2(byp_alu_rs1_data_e[8]), .Z(n1781) );
  HDINVD8 U2275 ( .A(ecl_shft_enshift_e_l), .Z(n2743) );
  HDINVD12 U2276 ( .A(byp_alu_rs2_data_e[4]), .Z(n3282) );
  HDINVDL U2277 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n228), .Z(
        n2467) );
  HDINVD1 U2278 ( .A(n2384), .Z(n2383) );
  HDNOR2D1 U2279 ( .A1(n3508), .A2(n3563), .Z(n2352) );
  HDNOR2D1 U2280 ( .A1(n3509), .A2(n3560), .Z(n2353) );
  HDNOR2M1D1 U2281 ( .A1(n2688), .A2(n3136), .Z(n2535) );
  HDINVD4 U2282 ( .A(n3569), .Z(n3487) );
  HDINVD8 U2283 ( .A(n3040), .Z(n2906) );
  HDNAN2D1 U2284 ( .A1(n2491), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n544), .Z(n2436) );
  HDBUFD8 U2285 ( .A(n3533), .Z(n2686) );
  HDINVD2 U2286 ( .A(n2675), .Z(n2015) );
  HDINVD4 U2287 ( .A(n3260), .Z(n3176) );
  HDINVBD2 U2288 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n140), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n571) );
  HDNOR2D4 U2289 ( .A1(n2725), .A2(ecl_shft_enshift_e_l), .Z(n3445) );
  HDINVD1 U2290 ( .A(byp_alu_rs2_data_e[27]), .Z(n2452) );
  HDINVD12 U2291 ( .A(ecl_alu_out_sel_logic_e_l), .Z(n2756) );
  HDINVD1 U2292 ( .A(byp_alu_rs1_data_e[38]), .Z(n3477) );
  HDINVD1 U2293 ( .A(byp_alu_rs1_data_e[26]), .Z(n2152) );
  HDINVD1 U2294 ( .A(byp_alu_rs1_data_e[17]), .Z(n1826) );
  HDINVD1 U2295 ( .A(byp_alu_rs2_data_e[62]), .Z(n2144) );
  HDINVD1 U2296 ( .A(byp_alu_rs2_data_e[49]), .Z(n2149) );
  HDINVD1 U2297 ( .A(byp_alu_rs2_data_e[53]), .Z(n1923) );
  HDINVD1 U2298 ( .A(ecl_alu_out_sel_shift_e_l), .Z(n1924) );
  HDINVD1 U2299 ( .A(byp_alu_rs2_data_e[34]), .Z(n1960) );
  HDINVD1 U2300 ( .A(byp_alu_rs1_data_e[28]), .Z(n2154) );
  HDINVD1 U2301 ( .A(byp_alu_rs1_data_e[35]), .Z(n3448) );
  HDNAN2M1D1 U2302 ( .A1(n2674), .A2(n2759), .Z(alu_byp_rd_data_e[0]) );
  HDOA222D1 U2303 ( .A1(n2923), .A2(n3561), .B1(n2881), .B2(n2702), .C1(n2905), 
        .C2(n3563), .Z(n2458) );
  HDOA22D1 U2304 ( .A1(n3326), .A2(n3576), .B1(n3325), .B2(n1783), .Z(n1933)
         );
  HDOA22D1 U2305 ( .A1(n3326), .A2(n3561), .B1(n3325), .B2(n1789), .Z(n1944)
         );
  HDOAI211D1 U2306 ( .A1(n3062), .A2(n3566), .B(n2723), .C(n1876), .Z(n2724)
         );
  HDINVD1 U2307 ( .A(n3308), .Z(n3164) );
  HDINVD4 U2308 ( .A(n2679), .Z(n2677) );
  HDINVD1 U2309 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n682), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n676) );
  HDNAN2D1 U2310 ( .A1(n2501), .A2(n2500), .Z(n2582) );
  HDOAI22D1 U2311 ( .A1(n2822), .A2(n1783), .B1(n2817), .B2(n3576), .Z(n2809)
         );
  HDOAI22D1 U2312 ( .A1(n2807), .A2(n1783), .B1(n2817), .B2(n3560), .Z(n2794)
         );
  HDOR2D1 U2313 ( .A1(n3369), .A2(n3576), .Z(n2082) );
  HDINVD2 U2314 ( .A(n3323), .Z(n3202) );
  HDINVD12 U2315 ( .A(n2977), .Z(n2908) );
  HDAOI22D1 U2316 ( .A1(n1975), .A2(n3192), .B1(n3191), .B2(
        byp_alu_rs1_data_e[28]), .Z(n3194) );
  HDNAN2M1D1 U2317 ( .A1(n2227), .A2(n1769), .Z(n2226) );
  HDAOI21D1 U2318 ( .A1(n3561), .A2(n3560), .B(n3575), .Z(n3577) );
  HDINVD1 U2319 ( .A(byp_alu_rs1_data_e[39]), .Z(n3486) );
  HDINVD1 U2320 ( .A(byp_alu_rs1_data_e[0]), .Z(n2670) );
  HDINVD1 U2321 ( .A(byp_alu_rs2_data_e[59]), .Z(n1829) );
  HDOA22M10D1 U2322 ( .A2(n3309), .A1(n1788), .B1(n3310), .B2(n3560), .Z(n1957) );
  HDAOI211D2 U2323 ( .A1(ecl_shft_shift4_e[2]), .A2(n3502), .B(n3456), .C(
        n3430), .Z(n3453) );
  HDAOI22D1 U2324 ( .A1(n2196), .A2(n2860), .B1(n2859), .B2(
        byp_alu_rs1_data_e[7]), .Z(n2862) );
  HDOAI22D1 U2325 ( .A1(n2977), .A2(n3383), .B1(n3498), .B2(n3040), .Z(n2925)
         );
  HDOAI22D1 U2326 ( .A1(n2977), .A2(n3394), .B1(n3505), .B2(n3040), .Z(n2943)
         );
  HDINVD1 U2327 ( .A(n3533), .Z(n1787) );
  HDNAN2D8 U2328 ( .A1(n2684), .A2(ecl_shft_shift4_e[3]), .Z(n3165) );
  HDNOR2D1 U2329 ( .A1(n2673), .A2(n2670), .Z(n2665) );
  HDINVBD2 U2330 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n95), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n93) );
  HDNAN2D1 U2331 ( .A1(n1767), .A2(n1862), .Z(n2521) );
  HDNAN2D1 U2332 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n996), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n848), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n613) );
  HDNAN2DL U2333 ( .A1(alu_addsub_rs2_data[31]), .A2(n1767), .Z(n3251) );
  HDNAN2M1D1 U2334 ( .A1(n1784), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n571), .Z(n2349) );
  HDINVBD20 U2335 ( .A(n1776), .Z(n1782) );
  HDAND2D1 U2336 ( .A1(n2138), .A2(byp_alu_rs1_data_e[30]), .Z(n2204) );
  HDNAN2D1 U2337 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n442), .A2(
        n2492), .Z(n2430) );
  HDINVD1 U2338 ( .A(n3431), .Z(n2883) );
  HDINVBD12 U2339 ( .A(n2688), .Z(n1789) );
  HDOR2D1 U2340 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_26_), .A2(
        byp_alu_rs1_data_e[58]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n569) );
  HDNAN2M1D1 U2341 ( .A1(n2310), .A2(n2027), .Z(n2026) );
  HDOAI22D1 U2342 ( .A1(n3300), .A2(n3561), .B1(n3299), .B2(n1789), .Z(n3274)
         );
  HDNOR2D1 U2343 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n738), .A2(
        n2112), .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n684) );
  HDOAI22D1 U2344 ( .A1(n3270), .A2(n3576), .B1(n3269), .B2(n1783), .Z(n3248)
         );
  HDOA22D1 U2345 ( .A1(n3415), .A2(n2702), .B1(n2590), .B2(n3533), .Z(n2461)
         );
  HDOR2D1 U2346 ( .A1(n3377), .A2(n3561), .Z(n2500) );
  HDOA22D1 U2347 ( .A1(n3377), .A2(n2702), .B1(n3376), .B2(n3533), .Z(n2048)
         );
  HDOA22D1 U2348 ( .A1(n3397), .A2(n3561), .B1(n3396), .B2(n1789), .Z(n2047)
         );
  HDNOR2M1D1 U2349 ( .A1(ecl_alu_out_sel_shift_e_l), .A2(n2565), .Z(n2562) );
  HDNOR2D1 U2350 ( .A1(n3326), .A2(n2702), .Z(n2069) );
  HDOA211D2 U2351 ( .A1(n3158), .A2(n2704), .B(n3102), .C(n3101), .Z(n3135) );
  HDOR2D1 U2352 ( .A1(n3299), .A2(n2686), .Z(n1940) );
  HDOA22D1 U2353 ( .A1(n3492), .A2(n3561), .B1(n2591), .B2(n1789), .Z(n1919)
         );
  HDAOI211D2 U2354 ( .A1(ecl_shft_shift4_e[3]), .A2(n3317), .B(n2237), .C(
        n2238), .Z(n3333) );
  HDINVD1 U2355 ( .A(n3487), .Z(n2126) );
  HDOR2D1 U2356 ( .A1(n3378), .A2(n2456), .Z(n2448) );
  HDAOI22D1 U2357 ( .A1(alu_addsub_rs2_data[13]), .A2(n2953), .B1(n2952), .B2(
        byp_alu_rs1_data_e[13]), .Z(n2955) );
  HDINVD1 U2358 ( .A(n3200), .Z(n3010) );
  HDNOR2D1 U2359 ( .A1(n3224), .A2(n2456), .Z(n3016) );
  HDINVBD2 U2360 ( .A(n3317), .Z(n3183) );
  HDOAI21M20D2 U2361 ( .A1(n3483), .A2(n2681), .B(n3095), .Z(n3308) );
  HDNOR2D1 U2362 ( .A1(n2672), .A2(n2135), .Z(n2664) );
  HDOAI21M20D1 U2363 ( .A1(n1782), .A2(n3008), .B(n3260), .Z(n3009) );
  HDNAN2D1 U2364 ( .A1(n2662), .A2(byp_alu_rs1_data_e[56]), .Z(n3497) );
  HDNAN2D1 U2365 ( .A1(n2690), .A2(byp_alu_rs1_data_e[21]), .Z(n2143) );
  HDNAN2D1 U2366 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n595), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n561), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n36) );
  HDOR2D1 U2367 ( .A1(n2290), .A2(ecl_alu_out_sel_sum_e_l), .Z(n2280) );
  HDINVD1 U2368 ( .A(n2255), .Z(n2271) );
  HDINVD1 U2369 ( .A(n1781), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n1002) );
  HDINVBD12 U2370 ( .A(n3549), .Z(n3576) );
  HDAND2D1 U2371 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n68), .A2(
        n2482), .Z(n2290) );
  HDNOR2D1 U2372 ( .A1(n2266), .A2(ecl_alu_out_sel_sum_e_l), .Z(n2255) );
  HDAND2D1 U2373 ( .A1(n2656), .A2(byp_alu_rs1_data_e[16]), .Z(n3265) );
  HDINVD1 U2374 ( .A(n1997), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n988) );
  HDINVD1 U2375 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n50), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n565) );
  HDOR2D1 U2376 ( .A1(alu_addsub_rs2_data[31]), .A2(byp_alu_rs1_data_e[31]), 
        .Z(n2496) );
  HDNOR2D2 U2377 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_24_), 
        .A2(byp_alu_rs1_data_e[56]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n140) );
  HDINVD16 U2378 ( .A(byp_alu_rs2_data_e[2]), .Z(n1797) );
  HDINVD1 U2379 ( .A(byp_alu_rs1_data_e[61]), .Z(n2289) );
  HDNOR2M1D2 U2380 ( .A1(n1959), .A2(n1952), .Z(n1949) );
  HDNAN2M1D1 U2381 ( .A1(ecl_alu_out_sel_shift_e_l), .A2(n2623), .Z(n2622) );
  HDOAI22D1 U2382 ( .A1(n3226), .A2(n3560), .B1(n3225), .B2(n3563), .Z(n2184)
         );
  HDOR2D1 U2383 ( .A1(n3300), .A2(n2702), .Z(n1939) );
  HDOA22D1 U2384 ( .A1(n3491), .A2(n3561), .B1(n3471), .B2(n3560), .Z(n1858)
         );
  HDOR2D1 U2385 ( .A1(n3376), .A2(n1789), .Z(n2501) );
  HDAOI211D2 U2386 ( .A1(ecl_shft_shift4_e[2]), .A2(n3323), .B(n3290), .C(
        n3289), .Z(n3309) );
  HDOA22D1 U2387 ( .A1(n3453), .A2(n3561), .B1(n3452), .B2(n1789), .Z(n1966)
         );
  HDOA22D1 U2388 ( .A1(n3451), .A2(n3560), .B1(n3450), .B2(n3563), .Z(n1964)
         );
  HDOA22D2 U2389 ( .A1(n3361), .A2(n3576), .B1(n2206), .B2(n1783), .Z(n1974)
         );
  HDOA22D1 U2390 ( .A1(n3433), .A2(n3560), .B1(n3432), .B2(n3563), .Z(n2460)
         );
  HDNAN2D1 U2391 ( .A1(n2760), .A2(ecl_shft_shift4_e[0]), .Z(n2763) );
  HDNOR2D1 U2392 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n395), .A2(
        n1790), .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n376) );
  HDAOI211D2 U2393 ( .A1(ecl_shft_shift4_e[3]), .A2(n3520), .B(n3410), .C(
        n3409), .Z(n3433) );
  HDAND2D2 U2394 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n366), .A2(
        n2375), .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n362) );
  HDAOI211D2 U2395 ( .A1(ecl_shft_shift4_e[3]), .A2(n3308), .B(n3306), .C(
        n3307), .Z(n3325) );
  HDAOI211D2 U2396 ( .A1(ecl_shft_shift4_e[0]), .A2(n3461), .B(n3351), .C(
        n3350), .Z(n3376) );
  HDNAN2D1 U2397 ( .A1(n2775), .A2(ecl_shft_shift4_e[0]), .Z(n2778) );
  HDAND3D1 U2398 ( .A1(n2442), .A2(n2443), .A3(n2444), .Z(n2437) );
  HDAOI22D1 U2399 ( .A1(alu_addsub_rs2_data[12]), .A2(n2937), .B1(n2936), .B2(
        byp_alu_rs1_data_e[12]), .Z(n2939) );
  HDAOI22D1 U2400 ( .A1(n2174), .A2(n2973), .B1(n2972), .B2(
        byp_alu_rs1_data_e[14]), .Z(n2975) );
  HDOR2D1 U2401 ( .A1(n2665), .A2(n2664), .Z(n2140) );
  HDAOI22D1 U2402 ( .A1(n1866), .A2(n3171), .B1(n3170), .B2(
        byp_alu_rs1_data_e[27]), .Z(n3173) );
  HDNAN2D1 U2403 ( .A1(n3569), .A2(ecl_shft_shift4_e[2]), .Z(n3523) );
  HDAOI22D1 U2404 ( .A1(n1978), .A2(n3233), .B1(n3232), .B2(
        byp_alu_rs1_data_e[30]), .Z(n3235) );
  HDAOI22D1 U2405 ( .A1(n1968), .A2(n3212), .B1(n3211), .B2(
        byp_alu_rs1_data_e[29]), .Z(n3214) );
  HDOA222D1 U2406 ( .A1(n1986), .A2(n2704), .B1(n3374), .B2(n2708), .C1(n3341), 
        .C2(n2710), .Z(n2577) );
  HDAOI22D1 U2407 ( .A1(n2136), .A2(n3277), .B1(n3276), .B2(
        byp_alu_rs1_data_e[32]), .Z(n3280) );
  HDOAI22D1 U2408 ( .A1(n2977), .A2(n3553), .B1(n3513), .B2(n3040), .Z(n2957)
         );
  HDAOI21D2 U2409 ( .A1(n2681), .A2(n3301), .B(n2327), .Z(n3240) );
  HDAND2D2 U2410 ( .A1(n3142), .A2(n2298), .Z(n3332) );
  HDOR2D1 U2411 ( .A1(n3416), .A2(n2704), .Z(n2449) );
  HDOA21D1 U2412 ( .A1(n2703), .A2(byp_alu_rs1_data_e[0]), .B(n1769), .Z(n2672) );
  HDINVD1 U2413 ( .A(n2436), .Z(n2435) );
  HDINVD1 U2414 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n688), .Z(
        n2112) );
  HDNOR2M1D1 U2415 ( .A1(n1785), .A2(n2291), .Z(n2281) );
  HDINVD1 U2416 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n561), .Z(
        n2195) );
  HDINVD1 U2417 ( .A(n2233), .Z(n2232) );
  HDOAI21M20D2 U2418 ( .A1(byp_alu_rs1_data_e[53]), .A2(n2745), .B(n2678), .Z(
        n3327) );
  HDNAN2D1 U2419 ( .A1(n2349), .A2(n1785), .Z(n2340) );
  HDINVD1 U2420 ( .A(n2290), .Z(n2291) );
  HDNAN2D1 U2421 ( .A1(n1767), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_29_), .Z(n2288) );
  HDINVD1 U2422 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n714), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n712) );
  HDNAN2D1 U2423 ( .A1(n1767), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_24_), .Z(n2348) );
  HDNAN2D1 U2424 ( .A1(n1767), .A2(n2183), .Z(n2425) );
  HDNAN2D1 U2425 ( .A1(n1767), .A2(n1980), .Z(n2405) );
  HDNAN2D1 U2426 ( .A1(n1767), .A2(n2161), .Z(n2641) );
  HDNAN2D1 U2427 ( .A1(alu_addsub_rs2_data[63]), .A2(n1767), .Z(n2257) );
  HDNAN2D1 U2428 ( .A1(n1767), .A2(n1999), .Z(n2541) );
  HDINVD1 U2429 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n777), .Z(
        n2357) );
  HDAND2D1 U2430 ( .A1(n2656), .A2(byp_alu_rs1_data_e[27]), .Z(n3375) );
  HDAND2D1 U2431 ( .A1(n2656), .A2(byp_alu_rs1_data_e[17]), .Z(n3288) );
  HDINVD1 U2432 ( .A(n2464), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n1006) );
  HDINVD1 U2433 ( .A(n2167), .Z(n2153) );
  HDNAN2D2 U2434 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_24_), 
        .A2(byp_alu_rs1_data_e[56]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n141) );
  HDNAN2D2 U2435 ( .A1(n2743), .A2(byp_alu_rs1_data_e[2]), .Z(n3436) );
  HDNAN2D1 U2436 ( .A1(n1731), .A2(byp_alu_rs1_data_e[16]), .Z(n1871) );
  HDNAN2D2 U2437 ( .A1(n2743), .A2(byp_alu_rs1_data_e[0]), .Z(n3422) );
  HDAND2D2 U2438 ( .A1(byp_alu_rs1_data_e[5]), .A2(n2743), .Z(n3464) );
  HDOA21D1 U2439 ( .A1(n2135), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n976), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n977), .Z(n2475) );
  HDNAN2D1 U2440 ( .A1(n2176), .A2(byp_alu_rs1_data_e[1]), .Z(n1872) );
  HDINVD1 U2441 ( .A(byp_alu_rs1_data_e[22]), .Z(n2586) );
  HDINVD1 U2442 ( .A(byp_alu_rs1_data_e[47]), .Z(n3568) );
  HDINVD1 U2443 ( .A(byp_alu_rs1_data_e[36]), .Z(n2248) );
  HDINVD8 U2444 ( .A(ecl_shft_extendbit_e), .Z(n3575) );
  HDINVD1 U2445 ( .A(byp_alu_rs1_data_e[49]), .Z(n2216) );
  HDOAI211D1 U2446 ( .A1(n2993), .A2(ecl_alu_out_sel_shift_e_l), .B(n2992), 
        .C(n2991), .Z(alu_byp_rd_data_e[15]) );
  HDOAI211D1 U2447 ( .A1(ecl_alu_out_sel_shift_e_l), .A2(n2880), .B(n2879), 
        .C(n2878), .Z(alu_byp_rd_data_e[8]) );
  HDOAI211D1 U2448 ( .A1(n2922), .A2(ecl_alu_out_sel_shift_e_l), .B(n2921), 
        .C(n2920), .Z(alu_byp_rd_data_e[11]) );
  HDOAI211D1 U2449 ( .A1(n2903), .A2(ecl_alu_out_sel_shift_e_l), .B(n2902), 
        .C(n2901), .Z(alu_byp_rd_data_e[10]) );
  HDOAI211D1 U2450 ( .A1(n3056), .A2(ecl_alu_out_sel_shift_e_l), .B(n3055), 
        .C(n3054), .Z(alu_byp_rd_data_e[19]) );
  HDOAI211D1 U2451 ( .A1(n2956), .A2(ecl_alu_out_sel_shift_e_l), .B(n2955), 
        .C(n2954), .Z(alu_byp_rd_data_e[13]) );
  HDOAI211D1 U2452 ( .A1(n2847), .A2(ecl_alu_out_sel_shift_e_l), .B(n2846), 
        .C(n2845), .Z(alu_byp_rd_data_e[6]) );
  HDOAI211D1 U2453 ( .A1(ecl_alu_out_sel_shift_e_l), .A2(n2940), .B(n2939), 
        .C(n2938), .Z(alu_byp_rd_data_e[12]) );
  HDOAI211D1 U2454 ( .A1(n2831), .A2(ecl_alu_out_sel_shift_e_l), .B(n2830), 
        .C(n2829), .Z(alu_byp_rd_data_e[5]) );
  HDNAN3D2 U2455 ( .A1(n2097), .A2(n2098), .A3(n2099), .Z(n2101) );
  HDOA22D1 U2456 ( .A1(n3572), .A2(n3563), .B1(n3573), .B2(n1783), .Z(n2614)
         );
  HDOA211D2 U2457 ( .A1(n2887), .A2(n2709), .B(n2763), .C(n2762), .Z(n2802) );
  HDNOR2D1 U2458 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n764), .A2(
        n2185), .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n749) );
  HDOA22D1 U2459 ( .A1(n3300), .A2(n3576), .B1(n3299), .B2(n1783), .Z(n1956)
         );
  HDOR2D1 U2460 ( .A1(n3342), .A2(n3563), .Z(n2074) );
  HDNOR2D1 U2461 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n738), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n725), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n723) );
  HDOA21M10D1 U2462 ( .A2(n3525), .A1(n2687), .B(n2646), .Z(n2648) );
  HDNOR2D2 U2463 ( .A1(n3222), .A2(n3221), .Z(n3292) );
  HDOA211D2 U2464 ( .A1(n2912), .A2(n2709), .B(n2791), .C(n2790), .Z(n2836) );
  HDOA211D2 U2465 ( .A1(n2892), .A2(n2707), .B(n2778), .C(n2777), .Z(n2817) );
  HDAOI211D2 U2466 ( .A1(ecl_shft_shift4_e[0]), .A2(n3554), .B(n3516), .C(
        n3517), .Z(n3534) );
  HDOAI21D1 U2467 ( .A1(n2459), .A2(n2476), .B(n1815), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n802) );
  HDAOI22D1 U2468 ( .A1(byp_alu_rs2_data_e[3]), .A2(n2683), .B1(
        alu_adder_out[3]), .B2(n1785), .Z(n2799) );
  HDAOI211D2 U2469 ( .A1(ecl_shft_shift4_e[2]), .A2(n3308), .B(n3244), .C(
        n3243), .Z(n3293) );
  HDAOI211D2 U2470 ( .A1(ecl_shft_shift4_e[3]), .A2(n3298), .B(n2328), .C(
        n2329), .Z(n2301) );
  HDOA21D1 U2471 ( .A1(n2419), .A2(n2414), .B(n2420), .Z(n2432) );
  HDAOI211D2 U2472 ( .A1(ecl_shft_shift4_e[2]), .A2(n3317), .B(n3268), .C(
        n3267), .Z(n3299) );
  HDOA22D1 U2473 ( .A1(n3296), .A2(n2456), .B1(n3328), .B2(n2704), .Z(n2004)
         );
  HDOA211D2 U2474 ( .A1(n3383), .A2(n1806), .B(n3382), .C(n3381), .Z(n2001) );
  HDNAN2D1 U2475 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n431), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n363), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n361) );
  HDAND2D1 U2476 ( .A1(n2435), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n561), .Z(n1995) );
  HDINVD1 U2477 ( .A(n2413), .Z(n2412) );
  HDNAN2D1 U2478 ( .A1(n2413), .A2(n1785), .Z(n2397) );
  HDAOI22D1 U2479 ( .A1(n2403), .A2(byp_alu_rs1_data_e[44]), .B1(n1980), .B2(
        n2404), .Z(n2401) );
  HDAOI22D1 U2480 ( .A1(byp_alu_rs1_data_e[52]), .A2(n1849), .B1(n1850), .B2(
        n1808), .Z(n1847) );
  HDAOI22D1 U2481 ( .A1(n2176), .A2(n2770), .B1(n2769), .B2(
        byp_alu_rs1_data_e[1]), .Z(n2771) );
  HDOAI21M20D2 U2482 ( .A1(n2138), .A2(byp_alu_rs1_data_e[33]), .B(n2504), .Z(
        n2583) );
  HDINVD1 U2483 ( .A(n2177), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n828) );
  HDOA21M10D1 U2484 ( .A2(n3414), .A1(n2662), .B(n2369), .Z(n3530) );
  HDAOI211D2 U2485 ( .A1(n2699), .A2(byp_alu_rs1_data_e[43]), .B(n2574), .C(
        n3375), .Z(n2124) );
  HDINVD12 U2486 ( .A(n2697), .Z(n2655) );
  HDAOI22D1 U2487 ( .A1(byp_alu_rs1_data_e[50]), .A2(n2518), .B1(n2519), .B2(
        n1861), .Z(n2516) );
  HDOA211D2 U2488 ( .A1(n3553), .A2(n2685), .B(n1730), .C(n2713), .Z(n2912) );
  HDNOR2D1 U2489 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n816), .A2(
        n2476), .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n801) );
  HDAOI22D1 U2490 ( .A1(n2193), .A2(n2844), .B1(n2843), .B2(
        byp_alu_rs1_data_e[6]), .Z(n2846) );
  HDINVBD2 U2491 ( .A(n2180), .Z(n2181) );
  HDINVD2 U2492 ( .A(n3407), .Z(n3239) );
  HDNAN2D1 U2493 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n688), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n662), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n660) );
  HDOAI21M20D2 U2494 ( .A1(n3124), .A2(n2681), .B(n3123), .Z(n3323) );
  HDNAN3D1 U2495 ( .A1(n1785), .A2(n2195), .A3(n2436), .Z(n2443) );
  HDAOI21D1 U2496 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n465), .A2(
        n2466), .B(n2142), .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n464)
         );
  HDINVBD4 U2497 ( .A(n1760), .Z(n3175) );
  HDNAN2D1 U2498 ( .A1(n1785), .A2(n2436), .Z(n2433) );
  HDNAN3D1 U2499 ( .A1(n1769), .A2(n2405), .A3(n2406), .Z(n2403) );
  HDNAN2D1 U2500 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n583), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n345), .Z(n2413) );
  HDNAN2D8 U2501 ( .A1(n1782), .A2(ecl_shft_shift4_e[2]), .Z(n3096) );
  HDINVD1 U2502 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n262), .Z(
        n2471) );
  HDOAI21M20D2 U2503 ( .A1(byp_alu_rs1_data_e[52]), .A2(n2745), .B(n2678), .Z(
        n3318) );
  HDINVD1 U2504 ( .A(n2465), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n906) );
  HDNAN2D1 U2505 ( .A1(n2233), .A2(n1785), .Z(n2219) );
  HDNAN2D1 U2506 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n1003), .A2(
        n1864), .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n620) );
  HDOAI21M20D2 U2507 ( .A1(byp_alu_rs1_data_e[54]), .A2(n2745), .B(n2676), .Z(
        n3336) );
  HDNAN2D1 U2508 ( .A1(n2313), .A2(n1785), .Z(n2310) );
  HDOR2D1 U2509 ( .A1(n1794), .A2(byp_alu_rs1_data_e[17]), .Z(n1793) );
  HDNAN2D1 U2510 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n980), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n643), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n597) );
  HDNAN2D1 U2511 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n953), .A2(
        n1810), .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n624) );
  HDNAN2D1 U2512 ( .A1(n2392), .A2(n1785), .Z(n2377) );
  HDNAN2D1 U2513 ( .A1(n2430), .A2(n1785), .Z(n2414) );
  HDNOR2D2 U2514 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n681), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n668), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n662) );
  HDINVD2 U2515 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n277), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n287) );
  HDINVD4 U2516 ( .A(n2202), .Z(n2700) );
  HDINVD2 U2517 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n72), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n82) );
  HDAND2D2 U2518 ( .A1(ifu_exu_invert_d), .A2(n1874), .Z(n1812) );
  HDNAN2D2 U2519 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I2_22_), 
        .A2(byp_alu_rs1_data_e[22]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n747) );
  HDINVD1 U2520 ( .A(n1808), .Z(n1853) );
  HDNAN2D2 U2521 ( .A1(n1886), .A2(byp_alu_rs1_data_e[19]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n778) );
  HDNAN2D2 U2522 ( .A1(n2147), .A2(byp_alu_rs1_data_e[18]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n799) );
  HDNAN2D2 U2523 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_3_), .A2(
        byp_alu_rs1_data_e[35]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n510) );
  HDOR2D1 U2524 ( .A1(n2130), .A2(byp_alu_rs1_data_e[24]), .Z(n2167) );
  HDNOR2D2 U2525 ( .A1(n1884), .A2(byp_alu_rs1_data_e[19]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n777) );
  HDNAN2D2 U2526 ( .A1(n2743), .A2(byp_alu_rs1_data_e[1]), .Z(n3431) );
  HDINVD1 U2527 ( .A(n1861), .Z(n2522) );
  HDNOR2D2 U2528 ( .A1(n2196), .A2(byp_alu_rs1_data_e[7]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n916) );
  HDNAN2D2 U2529 ( .A1(n1970), .A2(byp_alu_rs2_data_e[13]), .Z(n2166) );
  HDNAN2D2 U2530 ( .A1(ifu_exu_invert_d), .A2(n1816), .Z(n1817) );
  HDINVD2 U2531 ( .A(ecl_shft_shift4_e[2]), .Z(n2705) );
  HDOA31D2 U2532 ( .A1(ecl_shft_shift4_e[1]), .A2(ecl_shft_shift4_e[2]), .A3(
        ecl_shft_shift4_e[3]), .B(ecl_shft_extendbit_e), .Z(n3527) );
  HDINVD2 U2533 ( .A(byp_alu_rs1_data_e[3]), .Z(n2725) );
  HDEXOR2D2 U2534 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[31]), .Z(
        alu_addsub_rs2_data[31]) );
  HDNAN2D1 U2535 ( .A1(alu_addsub_rs2_data_1_), .A2(byp_alu_rs1_data_e[1]), 
        .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n969) );
  HDEXOR2D1 U2536 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[17]), .Z(
        alu_addsub_rs2_data[17]) );
  HDOR2D2 U2537 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n560), .A2(
        n2192), .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n531) );
  HDOA211D1 U2538 ( .A1(ecl_shft_op32_e), .A2(n2360), .B(byp_alu_rs2_data_e[4]), .C(n2743), .Z(n2656) );
  HDOAI22M20D1 U2539 ( .B1(n1928), .B2(ecl_alu_out_sel_shift_e_l), .A1(
        byp_alu_rs2_data_e[37]), .A2(n3579), .Z(n1927) );
  HDOA21M20D2 U2540 ( .A1(n2491), .A2(n2469), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n544), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n532) );
  HDOAI22M20D1 U2541 ( .B1(n1992), .B2(ecl_alu_out_sel_shift_e_l), .A1(n3579), 
        .A2(byp_alu_rs2_data_e[57]), .Z(n2373) );
  HDNOR2M1D1 U2542 ( .A1(ecl_shft_shift4_e[0]), .A2(n3493), .Z(n3494) );
  HDNOR3M1D1 U2543 ( .A1(ecl_shft_lshift_e_l), .A2(n1795), .A3(n3361), .Z(
        n2070) );
  HDOAI211D4 U2544 ( .A1(n2360), .A2(ecl_shft_op32_e), .B(n2743), .C(n3282), 
        .Z(n2202) );
  HDNOR2D1 U2545 ( .A1(n2272), .A2(n1737), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n963) );
  HDNAN2D2 U2546 ( .A1(n1746), .A2(byp_alu_rs2_data_e[2]), .Z(n1799) );
  HDNAN2D2 U2547 ( .A1(ifu_exu_invert_d), .A2(n1797), .Z(n1798) );
  HDEXOR2D1 U2548 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[1]), .Z(
        alu_addsub_rs2_data_1_) );
  HDEXOR2D1 U2549 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[0]), .Z(
        n1801) );
  HDOAI21M20D1 U2550 ( .A1(n1801), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n1010), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n977), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n975) );
  HDAOI21D1 U2551 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n963), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n975), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n964), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n962) );
  HDNAN2D1 U2552 ( .A1(n2333), .A2(byp_alu_rs1_data_e[3]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n960) );
  HDAOI21D1 U2553 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n945), .A2(
        n1881), .B(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n931), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n929) );
  HDNAN2D1 U2554 ( .A1(n1881), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n944), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n928) );
  HDOAI21D1 U2555 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n962), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n928), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n929), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n927) );
  HDAOI21D1 U2556 ( .A1(n2332), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n845), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n846), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n844) );
  HDOA21D2 U2557 ( .A1(n1888), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n843), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n844), .Z(n1802) );
  HDNOR2D1 U2558 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n883), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n843), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n841) );
  HDOA21M20D2 U2559 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n927), 
        .A2(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n841), .B(n1802), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n840) );
  HDEXOR2D1 U2560 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[22]), .Z(
        n1803) );
  HDOR2DL U2561 ( .A1(n2159), .A2(byp_alu_rs1_data_e[5]), .Z(n1805) );
  HDINVDL U2562 ( .A(n2697), .Z(n1806) );
  HDOA21D2 U2563 ( .A1(n3468), .A2(n3563), .B(n2094), .Z(n2099) );
  HDNAN2D2 U2564 ( .A1(ifu_exu_invert_d), .A2(n1983), .Z(n1984) );
  HDOA22D1 U2565 ( .A1(n3451), .A2(n3561), .B1(n3450), .B2(n1789), .Z(n2463)
         );
  HDEXOR2D1 U2566 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[43]), .Z(
        n1807) );
  HDNAN2DL U2567 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n992), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n799), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n609) );
  HDNOR2D2 U2568 ( .A1(byp_alu_rs1_data_e[0]), .A2(ecl_alu_cin_e), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n976) );
  HDNAN2D2 U2569 ( .A1(n1800), .A2(byp_alu_rs2_data_e[15]), .Z(n1818) );
  HDOA21D2 U2570 ( .A1(n3565), .A2(n1773), .B(n3242), .Z(n3374) );
  HDEXOR2D1 U2571 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[52]), .Z(
        n1809) );
  HDNAN2D2 U2572 ( .A1(n1971), .A2(byp_alu_rs2_data_e[18]), .Z(n1875) );
  HDNAN2D1 U2573 ( .A1(n2333), .A2(byp_alu_rs1_data_e[3]), .Z(n1810) );
  HDNOR2D2 U2574 ( .A1(n1812), .A2(n1813), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n798) );
  HDNAN2D2 U2575 ( .A1(n1875), .A2(n1811), .Z(n1813) );
  HDOA22D1 U2576 ( .A1(n3324), .A2(n2702), .B1(n2301), .B2(n3533), .Z(n1932)
         );
  HDOA22D1 U2577 ( .A1(n3324), .A2(n3561), .B1(n2301), .B2(n1789), .Z(n1955)
         );
  HDOA22D1 U2578 ( .A1(n3324), .A2(n3560), .B1(n2301), .B2(n3563), .Z(n1943)
         );
  HDNOR2D2 U2579 ( .A1(n1998), .A2(byp_alu_rs1_data_e[9]), .Z(n1814) );
  HDEXOR2D2 U2580 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[9]), .Z(
        n1998) );
  HDBUFDL U2581 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n804), .Z(
        n1815) );
  HDNAN2D2 U2582 ( .A1(n1817), .A2(n1818), .Z(alu_addsub_rs2_data_15_) );
  HDNAN2D2 U2583 ( .A1(alu_addsub_rs2_data_15_), .A2(byp_alu_rs1_data_e[15]), 
        .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n838) );
  HDOAI21D1 U2584 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n838), .A2(
        n2275), .B(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n825), .Z(n1821)
         );
  HDOA21M20D2 U2585 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n796), 
        .A2(n1821), .B(n1822), .Z(n1819) );
  HDOAI21D1 U2586 ( .A1(n1819), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n742), .B(n1893), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n737) );
  HDINVDL U2587 ( .A(n1819), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n793) );
  HDOAI21M20D1 U2588 ( .A1(n1843), .A2(n1785), .B(n1844), .Z(
        alu_byp_rd_data_e[59]) );
  HDOAI21D4 U2589 ( .A1(n1820), .A2(ecl_shft_op32_e), .B(byp_alu_rs2_data_e[4]), .Z(n2506) );
  HDOA21D1 U2590 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n804), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n798), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n799), .Z(n1822) );
  HDAOI21D1 U2591 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n663), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n640), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n641), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n639) );
  HDOA21D2 U2592 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n687), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n638), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n639), .Z(n1823) );
  HDOA21M20D2 U2593 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n636), 
        .A2(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n737), .B(n1823), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n635) );
  HDAOI22M10D1 U2594 ( .B1(n2653), .B2(byp_alu_rs1_data_e[33]), .A1(n1826), 
        .A2(n3550), .Z(n1825) );
  HDNAN2D1 U2595 ( .A1(n2700), .A2(byp_alu_rs1_data_e[49]), .Z(n1824) );
  HDOAI22D1 U2596 ( .A1(n3539), .A2(n2456), .B1(n2589), .B2(n2704), .Z(n1828)
         );
  HDNOR2D1 U2597 ( .A1(n2510), .A2(n2710), .Z(n1827) );
  HDAOI211D2 U2598 ( .A1(ecl_shft_shift4_e[2]), .A2(n3467), .B(n1827), .C(
        n1828), .Z(n3452) );
  HDOAI22DL U2599 ( .A1(n3564), .A2(n3561), .B1(n3545), .B2(n3560), .Z(n1837)
         );
  HDOAI22D1 U2600 ( .A1(n3526), .A2(n3576), .B1(n3519), .B2(n2702), .Z(n1836)
         );
  HDINVD1 U2601 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_27_), .Z(
        n1842) );
  HDNOR2D1 U2602 ( .A1(n1836), .A2(n1837), .Z(n1834) );
  HDNAN2D1 U2603 ( .A1(n1767), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_27_), .Z(n1841) );
  HDNAN2D1 U2604 ( .A1(n1772), .A2(n1842), .Z(n1840) );
  HDAOI21D1 U2605 ( .A1(n2481), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n125), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n126), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n124) );
  HDOAI22D1 U2606 ( .A1(n3534), .A2(n3563), .B1(n3544), .B2(n1789), .Z(n1833)
         );
  HDOAI211D1 U2607 ( .A1(n3518), .A2(n3533), .B(n1834), .C(n1835), .Z(n1832)
         );
  HDOAI21D1 U2608 ( .A1(n2703), .A2(byp_alu_rs1_data_e[59]), .B(n1769), .Z(
        n1839) );
  HDNAN3D1 U2609 ( .A1(n1769), .A2(n1840), .A3(n1841), .Z(n1838) );
  HDOR2D1 U2610 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n123), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n106), .Z(n1845) );
  HDAO21M20D1 U2611 ( .A1(n1832), .A2(n1833), .B(ecl_alu_out_sel_shift_e_l), 
        .Z(n1831) );
  HDAOI22D1 U2612 ( .A1(byp_alu_rs1_data_e[59]), .A2(n1838), .B1(n1839), .B2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_27_), .Z(n1830) );
  HDAOI21M20D2 U2613 ( .A1(n2012), .A2(n1845), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n105), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n103) );
  HDOA211D1 U2614 ( .A1(n2689), .A2(n1829), .B(n1830), .C(n1831), .Z(n1844) );
  HDEXOR2D2 U2615 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n103), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n9), .Z(n1843) );
  HDNAN2DL U2616 ( .A1(n1767), .A2(n1809), .Z(n1852) );
  HDNAN2D1 U2617 ( .A1(n1772), .A2(n1853), .Z(n1851) );
  HDOA22D1 U2618 ( .A1(n3469), .A2(n3576), .B1(n3453), .B2(n2702), .Z(n1859)
         );
  HDINVD1 U2619 ( .A(n3452), .Z(n1856) );
  HDOAI21D1 U2620 ( .A1(n2703), .A2(byp_alu_rs1_data_e[52]), .B(n1769), .Z(
        n1850) );
  HDNAN3D1 U2621 ( .A1(n1769), .A2(n1851), .A3(n1852), .Z(n1849) );
  HDOAI211D1 U2622 ( .A1(n3468), .A2(n1783), .B(n1858), .C(n1859), .Z(n1855)
         );
  HDAO22M10D1 U2623 ( .B1(n1856), .B2(n2687), .A2(n2688), .A1(n3490), .Z(n1854) );
  HDINVD1 U2624 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n226), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n224) );
  HDINVD1 U2625 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n225), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n223) );
  HDNAN2M1D1 U2626 ( .A1(n2689), .A2(byp_alu_rs2_data_e[52]), .Z(n1848) );
  HDNOR3M1D2 U2627 ( .A1(n1860), .A2(n1854), .A3(n1855), .Z(n1846) );
  HDAOI21D1 U2628 ( .A1(n2395), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n223), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n224), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n222) );
  HDOA211D1 U2629 ( .A1(n1846), .A2(ecl_alu_out_sel_shift_e_l), .B(n1847), .C(
        n1848), .Z(n1857) );
  HDOAI21M20D1 U2630 ( .A1(alu_adder_out_52_), .A2(n1785), .B(n1857), .Z(
        alu_byp_rd_data_e[52]) );
  HDEXOR2D1 U2631 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[50]), .Z(
        n1862) );
  HDEXOR2D1 U2632 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[50]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_18_) );
  HDOAI22D1 U2633 ( .A1(n2706), .A2(n3514), .B1(n2710), .B2(n3478), .Z(n3479)
         );
  HDNAN3D1 U2634 ( .A1(n1863), .A2(n2649), .A3(n2648), .Z(n2651) );
  HDOA22D1 U2635 ( .A1(n3534), .A2(n1783), .B1(n3573), .B2(n1789), .Z(n1863)
         );
  HDOA21M20D2 U2636 ( .A1(ecl_shft_shift4_e[1]), .A2(n3532), .B(n2550), .Z(
        n3573) );
  HDBUFD1 U2637 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n917), .Z(
        n1864) );
  HDNOR2D1 U2638 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n891), .A2(
        n1814), .Z(n1865) );
  HDNOR2D1 U2639 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n891), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n902), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n889) );
  HDEXOR2D1 U2640 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[27]), .Z(
        n1866) );
  HDNAN3D2 U2641 ( .A1(n2851), .A2(n3085), .A3(n2961), .Z(n3043) );
  HDAOI22DL U2642 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_22_), 
        .A2(n2225), .B1(n2226), .B2(byp_alu_rs1_data_e[54]), .Z(n2223) );
  HDMUX2DL U2643 ( .A0(n1772), .A1(n1767), .SL(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_22_), .Z(n2227) );
  HDEXNOR2D1 U2644 ( .A1(n3282), .A2(ifu_exu_invert_d), .Z(n2330) );
  HDINVD1 U2645 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n990), .Z(
        n1868) );
  HDEXOR2D1 U2646 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[42]), .Z(
        n1870) );
  HDNOR2D2 U2647 ( .A1(n3328), .A2(n2456), .Z(n3329) );
  HDOAI21M20D2 U2648 ( .A1(byp_alu_rs1_data_e[63]), .A2(n2745), .B(n2676), .Z(
        n3418) );
  HDOAI21M20D2 U2649 ( .A1(byp_alu_rs1_data_e[60]), .A2(n2745), .B(n2676), .Z(
        n3389) );
  HDOAI21M20D2 U2650 ( .A1(byp_alu_rs1_data_e[34]), .A2(n2745), .B(n2676), .Z(
        n3044) );
  HDOAI21M20D2 U2651 ( .A1(byp_alu_rs1_data_e[58]), .A2(n2745), .B(n2676), .Z(
        n3370) );
  HDOAI21M20D2 U2652 ( .A1(byp_alu_rs1_data_e[50]), .A2(n2745), .B(n2676), .Z(
        n3301) );
  HDEXOR2D1 U2653 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[7]), .Z(
        n2196) );
  HDNAN2D1 U2654 ( .A1(n2653), .A2(byp_alu_rs1_data_e[19]), .Z(n1876) );
  HDNAN2D1 U2655 ( .A1(n2653), .A2(byp_alu_rs1_data_e[19]), .Z(n3303) );
  HDNAN2DL U2656 ( .A1(n2832), .A2(ecl_shft_shift4_e[0]), .Z(n2835) );
  HDNOR2D1 U2657 ( .A1(n1927), .A2(n1929), .Z(n1926) );
  HDOAI211D2 U2658 ( .A1(n3331), .A2(n2654), .B(n2587), .C(n2507), .Z(n2508)
         );
  HDOAI22M10D1 U2659 ( .A1(n1766), .A2(n3471), .B1(n2702), .B2(n3451), .Z(
        n2095) );
  HDEXOR2D1 U2660 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[8]), .Z(
        n1878) );
  HDEXOR2D1 U2661 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[6]), .Z(
        n1879) );
  HDNAN2DL U2662 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n1002), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n914), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n619) );
  HDNAN2DL U2663 ( .A1(n1767), .A2(n1732), .Z(n2555) );
  HDEXOR2D1 U2664 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[6]), .Z(
        alu_addsub_rs2_data_6_) );
  HDNOR2D2 U2665 ( .A1(alu_addsub_rs2_data_6_), .A2(byp_alu_rs1_data_e[6]), 
        .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n932) );
  HDNOR2D2 U2666 ( .A1(n1879), .A2(byp_alu_rs1_data_e[6]), .Z(n2108) );
  HDNAN2DL U2667 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n994), .A2(
        n1871), .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n611) );
  HDNAN2D2 U2668 ( .A1(n1883), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n814), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n790) );
  HDAOI21D1 U2669 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n839), .A2(
        n1755), .B(n2474), .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n813)
         );
  HDNOR2D2 U2670 ( .A1(n2308), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n932), .Z(n1881) );
  HDNOR2D2 U2671 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n790), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n742), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n736) );
  HDINVD1 U2672 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n790), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n792) );
  HDNAN2D2 U2673 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n736), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n636), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n634) );
  HDOAI21DL U2674 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n840), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n634), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n635), .Z(n2479) );
  HDINVD1 U2675 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n796), .Z(
        n1882) );
  HDAOI22D1 U2676 ( .A1(n1885), .A2(n3053), .B1(n3052), .B2(
        byp_alu_rs1_data_e[19]), .Z(n3055) );
  HDEXOR2D1 U2677 ( .A1(byp_alu_rs2_data_e[19]), .A2(ifu_exu_invert_d), .Z(
        n1884) );
  HDEXOR2D1 U2678 ( .A1(byp_alu_rs2_data_e[19]), .A2(ifu_exu_invert_d), .Z(
        n1886) );
  HDEXOR2D1 U2679 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[8]), .Z(
        n1887) );
  HDNAN2D2 U2680 ( .A1(n1887), .A2(byp_alu_rs1_data_e[8]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n914) );
  HDAOI22DL U2681 ( .A1(n1887), .A2(n2877), .B1(n2876), .B2(
        byp_alu_rs1_data_e[8]), .Z(n2879) );
  HDOAI21D1 U2682 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n917), .A2(
        n1892), .B(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n914), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n908) );
  HDOAI21DL U2683 ( .A1(n1781), .A2(n1864), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n914), .Z(n2465) );
  HDOA21M20D2 U2684 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n908), 
        .A2(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n889), .B(n1891), .Z(
        n1888) );
  HDINVDL U2685 ( .A(n1888), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n886) );
  HDINVD2 U2686 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n737), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n739) );
  HDINVD4 U2687 ( .A(n2012), .Z(n1889) );
  HDAOI21D1 U2688 ( .A1(n1889), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n512), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n513), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n511) );
  HDAOI21D1 U2689 ( .A1(n1889), .A2(n1771), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n462), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n460) );
  HDNAN2D6 U2690 ( .A1(n2395), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n595), .Z(n2365) );
  HDAOI21D1 U2691 ( .A1(n1889), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n240), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n241), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n239) );
  HDAOI21D1 U2692 ( .A1(n2013), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n393), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n394), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n392) );
  HDAOI21D1 U2693 ( .A1(n1889), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n410), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n411), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n409) );
  HDINVBD4 U2694 ( .A(n2011), .Z(n1890) );
  HDAOI21D1 U2695 ( .A1(n1890), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n325), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n326), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n324) );
  HDAOI21D1 U2696 ( .A1(n1890), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n206), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n207), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n205) );
  HDAOI21D1 U2697 ( .A1(n1890), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n478), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n479), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n477) );
  HDAOI21D1 U2698 ( .A1(n1890), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n4), .B(n2481), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n290) );
  HDBUFBD4 U2699 ( .A(n1890), .Z(n2163) );
  HDOAI21M20D1 U2700 ( .A1(alu_adder_out_38_), .A2(n1785), .B(n2058), .Z(
        alu_byp_rd_data_e[38]) );
  HDOAI21M20D1 U2701 ( .A1(alu_adder_out_46_), .A2(n1785), .B(n1897), .Z(
        alu_byp_rd_data_e[46]) );
  HDOAI21M20D1 U2702 ( .A1(alu_adder_out_37_), .A2(n1785), .B(n1926), .Z(
        alu_byp_rd_data_e[37]) );
  HDOAI21M20D1 U2703 ( .A1(alu_adder_out_45_), .A2(n1785), .B(n1905), .Z(
        alu_byp_rd_data_e[45]) );
  HDOAI21M20D1 U2704 ( .A1(alu_adder_out_53_), .A2(n1785), .B(n1915), .Z(
        alu_byp_rd_data_e[53]) );
  HDOAI21M20D1 U2705 ( .A1(alu_adder_out_35_), .A2(n1785), .B(n1948), .Z(
        alu_byp_rd_data_e[35]) );
  HDOA21D1 U2706 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n891), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n903), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n892), .Z(n1891) );
  HDOAI21D1 U2707 ( .A1(n1997), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n752), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n747), .Z(n1894) );
  HDAOI21D1 U2708 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n767), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n744), .B(n1894), .Z(n1893)
         );
  HDNAN2D2 U2709 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n4), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n125), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n123) );
  HDOAI22D1 U2710 ( .A1(n3302), .A2(n2704), .B1(n3240), .B2(n2456), .Z(n1896)
         );
  HDNOR2D2 U2711 ( .A1(n3335), .A2(n2706), .Z(n1895) );
  HDAOI211D4 U2712 ( .A1(ecl_shft_shift4_e[3]), .A2(n3373), .B(n1895), .C(
        n1896), .Z(n3294) );
  HDOAI22M10D1 U2713 ( .A1(n1766), .A2(n3428), .B1(n1789), .B2(n3427), .Z(
        n1902) );
  HDOAI22D1 U2714 ( .A1(n3397), .A2(n2702), .B1(n3396), .B2(n2686), .Z(n1899)
         );
  HDOAI22D1 U2715 ( .A1(n3415), .A2(n3560), .B1(n2590), .B2(n3563), .Z(n1901)
         );
  HDINVD1 U2716 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n328), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n326) );
  HDINVD1 U2717 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n327), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n325) );
  HDNOR2D2 U2718 ( .A1(n1898), .A2(n1903), .Z(n1897) );
  HDMUXB2DL U2719 ( .A0(n1772), .A1(n1767), .SL(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_13_), .Z(n1912) );
  HDOAI22M10D1 U2720 ( .A1(n2503), .A2(n3395), .B1(n1914), .B2(n2686), .Z(
        n1911) );
  HDOAI22D1 U2721 ( .A1(n3397), .A2(n3576), .B1(n2114), .B2(n1783), .Z(n1908)
         );
  HDOAI22M10D1 U2722 ( .A1(n1766), .A2(n3415), .B1(n2590), .B2(n1789), .Z(
        n1910) );
  HDNOR2DL U2723 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n361), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n344), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n342) );
  HDNOR2D2 U2724 ( .A1(n1906), .A2(n1913), .Z(n1905) );
  HDOA22D2 U2725 ( .A1(n3471), .A2(n3576), .B1(n3470), .B2(n1783), .Z(n1918)
         );
  HDMUXB2DL U2726 ( .A0(n1772), .A1(n1767), .SL(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_21_), .Z(n1917) );
  HDNAN4D1 U2727 ( .A1(n1918), .A2(n1919), .A3(n1920), .A4(n1921), .Z(n1925)
         );
  HDNOR2D1 U2728 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n225), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n208), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n206) );
  HDAO22M10D1 U2729 ( .B1(n1925), .B2(n1924), .A2(n3579), .A1(n1923), .Z(n1916) );
  HDNOR2D2 U2730 ( .A1(n1922), .A2(n1916), .Z(n1915) );
  HDINVDL U2731 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n499), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n497) );
  HDAND4D1 U2732 ( .A1(n1930), .A2(n1931), .A3(n1932), .A4(n1933), .Z(n1928)
         );
  HDMUXB2DL U2733 ( .A0(n1772), .A1(n1767), .SL(n1945), .Z(n1938) );
  HDAOI21D1 U2734 ( .A1(n1938), .A2(n1769), .B(n3448), .Z(n1936) );
  HDOAI21D1 U2735 ( .A1(n2703), .A2(byp_alu_rs1_data_e[35]), .B(n1769), .Z(
        n1935) );
  HDOA22D1 U2736 ( .A1(n3310), .A2(n3576), .B1(n3309), .B2(n1783), .Z(n1942)
         );
  HDAND2D1 U2737 ( .A1(n1939), .A2(n1940), .Z(n1941) );
  HDOAI21DL U2738 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n532), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n514), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n515), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n513) );
  HDAOI21DL U2739 ( .A1(n1935), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_3_), .B(n1936), .Z(n1946) );
  HDAND4D1 U2740 ( .A1(n1941), .A2(n1942), .A3(n1943), .A4(n1944), .Z(n1937)
         );
  HDOA211D1 U2741 ( .A1(n1937), .A2(ecl_alu_out_sel_shift_e_l), .B(n1946), .C(
        n1947), .Z(n1948) );
  HDMUXB2DL U2742 ( .A0(n1772), .A1(n1767), .SL(n1958), .Z(n1953) );
  HDNAN4D1 U2743 ( .A1(n1956), .A2(n1957), .A3(n1954), .A4(n1955), .Z(n1961)
         );
  HDAOI21D1 U2744 ( .A1(n1953), .A2(n1769), .B(n3438), .Z(n1951) );
  HDOAI21D1 U2745 ( .A1(n2703), .A2(byp_alu_rs1_data_e[34]), .B(n1769), .Z(
        n1950) );
  HDINVD1 U2746 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n531), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n529) );
  HDAO22M20D1 U2747 ( .A1(n1960), .A2(n2689), .B1(n1961), .B2(n1924), .Z(n1952) );
  HDAOI21D1 U2748 ( .A1(n2157), .A2(n1950), .B(n1951), .Z(n1959) );
  HDAOI21D1 U2749 ( .A1(n2013), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n529), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n530), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n528) );
  HDOAI21M20D1 U2750 ( .A1(alu_adder_out_34_), .A2(n1785), .B(n1949), .Z(
        alu_byp_rd_data_e[34]) );
  HDOAI22D1 U2751 ( .A1(n3531), .A2(n2456), .B1(n2106), .B2(n2704), .Z(n1963)
         );
  HDAOI211D2 U2752 ( .A1(n3461), .A2(ecl_shft_shift4_e[3]), .B(n1962), .C(
        n1963), .Z(n3490) );
  HDAOI22D1 U2753 ( .A1(n2683), .A2(byp_alu_rs2_data_e[19]), .B1(
        alu_adder_out[19]), .B2(n1785), .Z(n3054) );
  HDOA22D1 U2754 ( .A1(n3433), .A2(n3576), .B1(n3432), .B2(n1783), .Z(n1965)
         );
  HDAND4D1 U2755 ( .A1(n2009), .A2(n1964), .A3(n1965), .A4(n1966), .Z(n2214)
         );
  HDEXOR2D1 U2756 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[37]), .Z(
        n1967) );
  HDEXOR2D1 U2757 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[29]), .Z(
        n1968) );
  HDNAN3D2 U2758 ( .A1(n2036), .A2(n2037), .A3(n2038), .Z(n2032) );
  HDOA211D2 U2759 ( .A1(n3394), .A2(n2696), .B(n2339), .C(n3393), .Z(n2589) );
  HDNAN2D2 U2760 ( .A1(n1973), .A2(n1974), .Z(n1972) );
  HDOA22D1 U2761 ( .A1(n3369), .A2(n3560), .B1(n3368), .B2(n3563), .Z(n1973)
         );
  HDEXOR2D1 U2762 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[28]), .Z(
        n1975) );
  HDINVD1 U2763 ( .A(n1743), .Z(n2668) );
  HDOAI22D1 U2764 ( .A1(n3518), .A2(n1789), .B1(n3500), .B2(n1783), .Z(n2351)
         );
  HDOAI22M10D1 U2765 ( .A1(byp_alu_rs2_data_e[40]), .A2(n2689), .B1(n2580), 
        .B2(ecl_alu_out_sel_shift_e_l), .Z(n2579) );
  HDINVDL U2766 ( .A(n1748), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n990) );
  HDEXOR2D1 U2767 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[48]), .Z(
        n1977) );
  HDEXOR2D1 U2768 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[48]), .Z(
        n2451) );
  HDEXOR2D1 U2769 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[30]), .Z(
        n1978) );
  HDINVBD4 U2770 ( .A(n1768), .Z(n2699) );
  HDAOI211D4 U2771 ( .A1(ecl_shft_shift4_e[1]), .A2(n3367), .B(n3330), .C(
        n3329), .Z(n3361) );
  HDINVD2 U2772 ( .A(n1870), .Z(n2396) );
  HDEXOR2D1 U2773 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[44]), .Z(
        n1981) );
  HDEXOR2D1 U2774 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[44]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_12_) );
  HDNOR2D1 U2775 ( .A1(n2158), .A2(ecl_shft_op32_e), .Z(n1982) );
  HDNOR2D6 U2776 ( .A1(n2470), .A2(ecl_shft_enshift_e_l), .Z(n3550) );
  HDOAI21D1 U2777 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n430), .A2(
        n2122), .B(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n298), .Z(n2481)
         );
  HDNOR2D1 U2778 ( .A1(n1744), .A2(n3438), .Z(n3439) );
  HDAND2D1 U2779 ( .A1(n3571), .A2(n2688), .Z(n2613) );
  HDOR2D2 U2780 ( .A1(alu_addsub_rs2_data[33]), .A2(byp_alu_rs1_data_e[33]), 
        .Z(n2491) );
  HDNAN2D1 U2781 ( .A1(n2832), .A2(ecl_shft_shift4_e[2]), .Z(n2747) );
  HDNAN2D2 U2782 ( .A1(n1747), .A2(byp_alu_rs2_data_e[16]), .Z(n1985) );
  HDNAN2D2 U2783 ( .A1(n1984), .A2(n1985), .Z(alu_addsub_rs2_data[16]) );
  HDINVD4 U2784 ( .A(n2202), .Z(n2203) );
  HDOA211D1 U2785 ( .A1(n3305), .A2(n2694), .B(n3304), .C(n1876), .Z(n1986) );
  HDOAI22D1 U2786 ( .A1(n3519), .A2(n3560), .B1(n3518), .B2(n3563), .Z(n1987)
         );
  HDOAI22D1 U2787 ( .A1(n3501), .A2(n2702), .B1(n3500), .B2(n3533), .Z(n1988)
         );
  HDOR2D1 U2788 ( .A1(n1987), .A2(n1988), .Z(n1989) );
  HDOAI22D1 U2789 ( .A1(n3509), .A2(n3576), .B1(n3508), .B2(n1783), .Z(n1990)
         );
  HDOAI22D1 U2790 ( .A1(n3526), .A2(n3561), .B1(n3525), .B2(n1789), .Z(n1991)
         );
  HDNOR3D2 U2791 ( .A1(n1989), .A2(n1990), .A3(n1991), .Z(n1992) );
  HDOA21D2 U2792 ( .A1(n3320), .A2(n2696), .B(n2511), .Z(n1993) );
  HDAND2D2 U2793 ( .A1(n1993), .A2(n2509), .Z(n2510) );
  HDNOR2D1 U2794 ( .A1(n2510), .A2(n2704), .Z(n3360) );
  HDAOI211D2 U2795 ( .A1(n3449), .A2(ecl_shft_shift4_e[2]), .B(n2208), .C(
        n2209), .Z(n1994) );
  HDAOI211D2 U2796 ( .A1(n3449), .A2(ecl_shft_shift4_e[2]), .B(n2208), .C(
        n2209), .Z(n3432) );
  HDNAN3D2 U2797 ( .A1(n2365), .A2(n1785), .A3(n1995), .Z(n2366) );
  HDNOR2D2 U2798 ( .A1(n3015), .A2(n3014), .Z(n3224) );
  HDNOR2D2 U2799 ( .A1(n2654), .A2(n3521), .Z(n2574) );
  HDNAN2D2 U2800 ( .A1(n2743), .A2(byp_alu_rs1_data_e[11]), .Z(n3521) );
  HDNOR2D1 U2801 ( .A1(n3559), .A2(n2704), .Z(n3480) );
  HDINVD20 U2802 ( .A(ecl_shft_extend32bit_e_l), .Z(n2712) );
  HDOA211D1 U2803 ( .A1(n3383), .A2(n2694), .B(n3382), .C(n3381), .Z(n3499) );
  HDEXOR2D1 U2804 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[1]), .Z(
        n1996) );
  HDAOI211D2 U2805 ( .A1(ecl_shft_shift4_e[2]), .A2(n3373), .B(n2306), .C(
        n2307), .Z(n3326) );
  HDINVDL U2806 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n663), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n665) );
  HDINVD2 U2807 ( .A(n1778), .Z(n2105) );
  HDNOR2D2 U2808 ( .A1(n1803), .A2(byp_alu_rs1_data_e[22]), .Z(n1997) );
  HDNAN2D1 U2809 ( .A1(n2656), .A2(byp_alu_rs1_data_e[32]), .Z(n2368) );
  HDINVBD4 U2810 ( .A(n2695), .Z(n2696) );
  HDAOI211D2 U2811 ( .A1(n2701), .A2(byp_alu_rs1_data_e[50]), .B(n3440), .C(
        n3439), .Z(n2002) );
  HDAOI211D1 U2812 ( .A1(n2701), .A2(byp_alu_rs1_data_e[50]), .B(n3440), .C(
        n3439), .Z(n3559) );
  HDNOR2D1 U2813 ( .A1(n3478), .A2(n2456), .Z(n2363) );
  HDOR2D1 U2814 ( .A1(n3399), .A2(n2710), .Z(n2003) );
  HDOAI211D2 U2815 ( .A1(n3218), .A2(n2675), .B(n3260), .C(n3217), .Z(n3367)
         );
  HDAOI21M20D2 U2816 ( .A1(n2299), .A2(n3436), .B(n3297), .Z(n2362) );
  HDOAI22D2 U2817 ( .A1(n3179), .A2(n2704), .B1(n3111), .B2(n2456), .Z(n3116)
         );
  HDOA22DL U2818 ( .A1(n3240), .A2(n2709), .B1(n3302), .B2(n2710), .Z(n3101)
         );
  HDINVD4 U2819 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n297), .Z(
        n2121) );
  HDNAN2D2 U2820 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n299), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n363), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n297) );
  HDNOR2D1 U2821 ( .A1(n2589), .A2(n2706), .Z(n2618) );
  HDEXOR2D1 U2822 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[25]), .Z(
        n2006) );
  HDOA21M10D2 U2823 ( .A2(n3414), .A1(n2662), .B(n2369), .Z(n2106) );
  HDINVD2 U2824 ( .A(n3536), .Z(n2008) );
  HDOAI22D1 U2825 ( .A1(n2928), .A2(n2710), .B1(n2804), .B2(n2704), .Z(n2731)
         );
  HDOA22D2 U2826 ( .A1(n3428), .A2(n2702), .B1(n3427), .B2(n3533), .Z(n2009)
         );
  HDNAN2D2 U2827 ( .A1(byp_alu_rs1_data_e[25]), .A2(n2690), .Z(n3356) );
  HDOAI211D1 U2828 ( .A1(n3505), .A2(n2685), .B(n3356), .C(n2746), .Z(n2832)
         );
  HDOAI211D1 U2829 ( .A1(n3505), .A2(n2696), .B(n3357), .C(n3356), .Z(n3467)
         );
  HDNOR2D2 U2830 ( .A1(n1809), .A2(byp_alu_rs1_data_e[52]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n208) );
  HDAOI21M20D2 U2831 ( .A1(n3376), .A2(n3563), .B(n2080), .Z(n2079) );
  HDAOI211D2 U2832 ( .A1(ecl_shft_shift4_e[3]), .A2(n3457), .B(n2019), .C(
        n2020), .Z(n3377) );
  HDOAI22D2 U2833 ( .A1(n3257), .A2(n2708), .B1(n3178), .B2(n2710), .Z(n3115)
         );
  HDAOI211D4 U2834 ( .A1(ecl_shft_shift4_e[0]), .A2(n3314), .B(n3313), .C(
        n3312), .Z(n3334) );
  HDINVDL U2835 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n962), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n961) );
  HDINVD1 U2836 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n927), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n926) );
  HDINVBD8 U2837 ( .A(n1724), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n839) );
  HDOAI21M20D2 U2838 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n633), 
        .A2(n2496), .B(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n632), .Z(
        n2010) );
  HDINVBD4 U2839 ( .A(n2010), .Z(n2011) );
  HDINVBD2 U2840 ( .A(n2010), .Z(n2012) );
  HDINVD4 U2841 ( .A(n2011), .Z(n2013) );
  HDAOI21M10D1 U2842 ( .A1(n2011), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n257), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n258), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n256) );
  HDINVD2 U2843 ( .A(n2011), .Z(n2395) );
  HDNOR2D2 U2844 ( .A1(n2012), .A2(n2150), .Z(n2497) );
  HDAOI21D1 U2845 ( .A1(n2013), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n376), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n377), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n375) );
  HDAOI21D1 U2846 ( .A1(n2013), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n121), .B(n2129), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n120) );
  HDBUFBD4 U2847 ( .A(n2013), .Z(n2190) );
  HDAOI21D1 U2848 ( .A1(n1889), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n499), .B(n2466), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n494) );
  HDAOI21D1 U2849 ( .A1(n2013), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n431), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n432), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n426) );
  HDOAI21M20D1 U2850 ( .A1(alu_adder_out_42_), .A2(n1785), .B(n2049), .Z(
        alu_byp_rd_data_e[42]) );
  HDOAI21M20D1 U2851 ( .A1(alu_adder_out_41_), .A2(n1785), .B(n2075), .Z(
        alu_byp_rd_data_e[41]) );
  HDOAI21M20D1 U2852 ( .A1(alu_adder_out_51_), .A2(n1785), .B(n2103), .Z(
        alu_byp_rd_data_e[51]) );
  HDAOI211D4 U2853 ( .A1(n3120), .A2(n1782), .B(n3176), .C(n2014), .Z(n3319)
         );
  HDAND2D1 U2854 ( .A1(n1756), .A2(n2015), .Z(n2014) );
  HDNOR2D2 U2855 ( .A1(n3319), .A2(n2456), .Z(n2018) );
  HDOAI22D1 U2856 ( .A1(n3429), .A2(n2710), .B1(n3390), .B2(n2707), .Z(n2017)
         );
  HDAOI211D4 U2857 ( .A1(ecl_shft_shift4_e[1]), .A2(n3354), .B(n2017), .C(
        n2018), .Z(n3343) );
  HDOAI22D1 U2858 ( .A1(n3378), .A2(n2704), .B1(n3345), .B2(n2456), .Z(n2020)
         );
  HDNOR2D1 U2859 ( .A1(n3416), .A2(n2706), .Z(n2019) );
  HDAOI211D2 U2860 ( .A1(n3449), .A2(ecl_shft_shift4_e[1]), .B(n2576), .C(
        n2575), .Z(n3396) );
  HDOA21DL U2861 ( .A1(n2467), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n195), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n196), .Z(n2022) );
  HDOA21M20D2 U2862 ( .A1(n1754), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n193), .B(n2022), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n192) );
  HDOA21D2 U2863 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n192), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n174), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n175), .Z(n2311) );
  HDOAI222D1 U2864 ( .A1(n3501), .A2(n3560), .B1(n3492), .B2(n3576), .C1(n3509), .C2(n3561), .Z(n2035) );
  HDOR2D1 U2865 ( .A1(n2591), .A2(n1783), .Z(n2038) );
  HDOR2D1 U2866 ( .A1(n3491), .A2(n2702), .Z(n2037) );
  HDNOR2M1D1 U2867 ( .A1(byp_alu_rs2_data_e[55]), .A2(n2689), .Z(n2030) );
  HDOAI21D1 U2868 ( .A1(n2703), .A2(byp_alu_rs1_data_e[55]), .B(n1769), .Z(
        n2028) );
  HDAOI211D1 U2869 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_23_), 
        .A2(n2028), .B(n2029), .C(n2030), .Z(n2025) );
  HDOA22D1 U2870 ( .A1(n2031), .A2(ecl_alu_out_sel_shift_e_l), .B1(n2312), 
        .B2(n2310), .Z(n2023) );
  HDNAN4D1 U2871 ( .A1(n2023), .A2(n2024), .A3(n2025), .A4(n2026), .Z(
        alu_byp_rd_data_e[55]) );
  HDNAN2D1 U2872 ( .A1(n1767), .A2(n1807), .Z(n2044) );
  HDNAN2D1 U2873 ( .A1(n1772), .A2(n2588), .Z(n2043) );
  HDOA22D1 U2874 ( .A1(n3388), .A2(n3576), .B1(n3387), .B2(n1783), .Z(n2046)
         );
  HDOA22D1 U2875 ( .A1(n3395), .A2(n3560), .B1(n2359), .B2(n3563), .Z(n2045)
         );
  HDNAN2M1D1 U2876 ( .A1(n2689), .A2(byp_alu_rs2_data_e[43]), .Z(n2042) );
  HDAND4D1 U2877 ( .A1(n2045), .A2(n2047), .A3(n2046), .A4(n2048), .Z(n2040)
         );
  HDOA211D1 U2878 ( .A1(n2040), .A2(ecl_alu_out_sel_shift_e_l), .B(n2041), .C(
        n2042), .Z(n2039) );
  HDOAI21M20D1 U2879 ( .A1(alu_adder_out_43_), .A2(n1785), .B(n2039), .Z(
        alu_byp_rd_data_e[43]) );
  HDNAN2DL U2880 ( .A1(n1767), .A2(n1870), .Z(n2054) );
  HDNAN2DL U2881 ( .A1(n1772), .A2(n2396), .Z(n2053) );
  HDOR2D1 U2882 ( .A1(n3395), .A2(n3561), .Z(n2057) );
  HDOAI211D1 U2883 ( .A1(n3376), .A2(n1783), .B(n2056), .C(n2057), .Z(n2055)
         );
  HDINVD1 U2884 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n396), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n394) );
  HDINVD1 U2885 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n395), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n393) );
  HDNAN2M1D1 U2886 ( .A1(n2689), .A2(byp_alu_rs2_data_e[42]), .Z(n2052) );
  HDOA211D1 U2887 ( .A1(n2050), .A2(ecl_alu_out_sel_shift_e_l), .B(n2051), .C(
        n2052), .Z(n2049) );
  HDINVDL U2888 ( .A(alu_addsub_rs2_data[38]), .Z(n2066) );
  HDNAN2DL U2889 ( .A1(n1767), .A2(alu_addsub_rs2_data[38]), .Z(n2065) );
  HDNAN2D1 U2890 ( .A1(n1772), .A2(n2066), .Z(n2064) );
  HDNOR2D1 U2891 ( .A1(n2206), .A2(n1789), .Z(n2071) );
  HDNAN3D1 U2892 ( .A1(n1769), .A2(n2064), .A3(n2065), .Z(n2063) );
  HDOAI21D1 U2893 ( .A1(n2703), .A2(byp_alu_rs1_data_e[38]), .B(n1769), .Z(
        n2062) );
  HDNAN2D2 U2894 ( .A1(n2073), .A2(n2074), .Z(n2072) );
  HDOR3D1 U2895 ( .A1(n2069), .A2(n2070), .A3(n2071), .Z(n2068) );
  HDINVD1 U2896 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n464), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n462) );
  HDNAN2M1D1 U2897 ( .A1(n2689), .A2(byp_alu_rs2_data_e[38]), .Z(n2061) );
  HDAOI22M10DL U2898 ( .B1(n2062), .B2(alu_addsub_rs2_data[38]), .A1(n3477), 
        .A2(n2063), .Z(n2060) );
  HDNOR3D2 U2899 ( .A1(n2068), .A2(n2072), .A3(n2067), .Z(n2059) );
  HDNAN2DL U2900 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n589), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n447), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n30) );
  HDOA211D1 U2901 ( .A1(n2059), .A2(ecl_alu_out_sel_shift_e_l), .B(n2060), .C(
        n2061), .Z(n2058) );
  HDNAN2D1 U2902 ( .A1(n1767), .A2(n2187), .Z(n2077) );
  HDINVDL U2903 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n430), .Z(
        n2088) );
  HDOAI22M10D1 U2904 ( .A1(n1787), .A2(n2206), .B1(n3377), .B2(n3560), .Z(
        n2080) );
  HDNAN3D2 U2905 ( .A1(n2082), .A2(n2083), .A3(n2084), .Z(n2081) );
  HDAOI21M20D2 U2906 ( .A1(n3368), .A2(n1783), .B(n2081), .Z(n2078) );
  HDOAI21DL U2907 ( .A1(n2089), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n412), .B(n2447), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n411) );
  HDNOR2DL U2908 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n429), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n412), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n410) );
  HDOA211D1 U2909 ( .A1(n3387), .A2(n1789), .B(n2078), .C(n2079), .Z(n2086) );
  HDOA211D1 U2910 ( .A1(n2086), .A2(ecl_alu_out_sel_shift_e_l), .B(n2085), .C(
        n2087), .Z(n2075) );
  HDOAI22D1 U2911 ( .A1(n3469), .A2(n3560), .B1(n3453), .B2(n3576), .Z(n2096)
         );
  HDNAN2D1 U2912 ( .A1(n1767), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_19_), .Z(n2093) );
  HDNOR2D2 U2913 ( .A1(n2096), .A2(n2095), .Z(n2094) );
  HDOAI21D1 U2914 ( .A1(n2703), .A2(byp_alu_rs1_data_e[51]), .B(n1769), .Z(
        n2091) );
  HDNAN3D1 U2915 ( .A1(n1769), .A2(n2092), .A3(n2093), .Z(n2090) );
  HDOA22D4 U2916 ( .A1(n3452), .A2(n1783), .B1(n3450), .B2(n3533), .Z(n2098)
         );
  HDNOR2D1 U2917 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n259), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n242), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n240) );
  HDAO22DL U2918 ( .A1(byp_alu_rs1_data_e[51]), .A2(n2090), .B1(n2091), .B2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_19_), .Z(n2102) );
  HDAOI211D1 U2919 ( .A1(n2101), .A2(n1924), .B(n2102), .C(n2100), .Z(n2103)
         );
  HDEXOR2D1 U2920 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[46]), .Z(
        n2104) );
  HDAOI22D1 U2921 ( .A1(n2697), .A2(n3088), .B1(n3536), .B2(n3327), .Z(n2740)
         );
  HDINVDL U2922 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n642), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n980) );
  HDINVDL U2923 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n651), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n981) );
  HDAOI22DL U2924 ( .A1(n2006), .A2(n3131), .B1(n3130), .B2(
        byp_alu_rs1_data_e[25]), .Z(n3133) );
  HDOAI211D1 U2925 ( .A1(n3498), .A2(n2654), .B(n3348), .C(n3347), .Z(n3461)
         );
  HDOAI22M10D1 U2926 ( .A1(n2786), .A2(n2693), .B1(n3436), .B2(n3566), .Z(
        n3440) );
  HDAOI211D2 U2927 ( .A1(ecl_shft_shift4_e[1]), .A2(n3314), .B(n3263), .C(
        n3262), .Z(n3300) );
  HDNAN2D2 U2928 ( .A1(n2107), .A2(n3446), .Z(n3569) );
  HDNAN2D1 U2929 ( .A1(n3550), .A2(byp_alu_rs1_data_e[19]), .Z(n3447) );
  HDEXOR2D1 U2930 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[23]), .Z(
        n2111) );
  HDEXOR2D2 U2931 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[23]), .Z(
        n2110) );
  HDNOR2D2 U2932 ( .A1(n3425), .A2(n2667), .Z(n3426) );
  HDAOI21D1 U2933 ( .A1(n3336), .A2(n2304), .B(n3176), .Z(n2305) );
  HDOAI22M10DL U2934 ( .A1(n1788), .A2(n3204), .B1(n3205), .B2(n3560), .Z(
        n3166) );
  HDOAI211D1 U2935 ( .A1(ecl_alu_out_sel_shift_e_l), .A2(n2317), .B(n2318), 
        .C(n2319), .Z(alu_byp_rd_data_e[22]) );
  HDAOI21D2 U2936 ( .A1(n2682), .A2(n3327), .B(n3089), .Z(n3296) );
  HDAOI22M10D1 U2937 ( .B1(n3536), .B2(n3398), .A1(n2655), .A2(n3216), .Z(
        n2742) );
  HDINVD1 U2938 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n686), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n688) );
  HDAO22M10D1 U2939 ( .B1(byp_alu_rs2_data_e[48]), .B2(n3579), .A2(n2113), 
        .A1(ecl_alu_out_sel_shift_e_l), .Z(n3425) );
  HDNAN4D1 U2940 ( .A1(n2460), .A2(n2461), .A3(n2462), .A4(n2463), .Z(n2113)
         );
  HDAOI211D2 U2941 ( .A1(n3532), .A2(ecl_shft_shift4_e[0]), .B(n2370), .C(
        n2371), .Z(n3518) );
  HDOAI211D1 U2942 ( .A1(n2863), .A2(ecl_alu_out_sel_shift_e_l), .B(n2862), 
        .C(n2861), .Z(alu_byp_rd_data_e[7]) );
  HDINVDL U2943 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n446), .Z(
        n2431) );
  HDAOI211D2 U2944 ( .A1(n3449), .A2(ecl_shft_shift4_e[1]), .B(n2576), .C(
        n2575), .Z(n2114) );
  HDINVD2 U2945 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n272), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n270) );
  HDNOR2D1 U2946 ( .A1(n3116), .A2(n3115), .Z(n2115) );
  HDNAN2DL U2947 ( .A1(n3550), .A2(byp_alu_rs1_data_e[23]), .Z(n3485) );
  HDAOI22DL U2948 ( .A1(n3550), .A2(byp_alu_rs1_data_e[29]), .B1(n2690), .B2(
        byp_alu_rs1_data_e[45]), .Z(n3538) );
  HDAND2DL U2949 ( .A1(n3550), .A2(byp_alu_rs1_data_e[28]), .Z(n2548) );
  HDINVDL U2950 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n707), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n985) );
  HDAOI211D1 U2951 ( .A1(byp_alu_rs1_data_e[32]), .A2(n2662), .B(n3265), .C(
        n3266), .Z(n2661) );
  HDEXOR2D1 U2952 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[26]), .Z(
        n2116) );
  HDINVD2 U2953 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n162), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n160) );
  HDAO21D2 U2954 ( .A1(n2508), .A2(ecl_shft_shift4_e[1]), .B(n2363), .Z(n2358)
         );
  HDINVD1 U2955 ( .A(n2118), .Z(n2119) );
  HDNAN2M1DL U2956 ( .A1(n1981), .A2(n1772), .Z(n2406) );
  HDNOR2D6 U2957 ( .A1(n3450), .A2(n1783), .Z(n2524) );
  HDAOI22M10D1 U2958 ( .B1(ecl_shft_shift4_e[3]), .B2(n3011), .A1(n2708), .A2(
        n2946), .Z(n2820) );
  HDEXOR2D1 U2959 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[40]), .Z(
        n2120) );
  HDOAI22DL U2960 ( .A1(n3564), .A2(n3576), .B1(n3545), .B2(n2702), .Z(n2296)
         );
  HDNOR2DL U2961 ( .A1(n3564), .A2(n2702), .Z(n2617) );
  HDOAI22M10D2 U2962 ( .A1(n3177), .A2(n2109), .B1(n3175), .B2(n2654), .Z(
        n2927) );
  HDNAN2D1 U2963 ( .A1(n2684), .A2(n3258), .Z(n3259) );
  HDOAI21M20D2 U2964 ( .A1(byp_alu_rs1_data_e[42]), .A2(n2745), .B(n2677), .Z(
        n3159) );
  HDOAI22M10D1 U2965 ( .A1(ecl_shft_shift4_e[3]), .A2(n3416), .B1(n3378), .B2(
        n2708), .Z(n3313) );
  HDOAI21M20D2 U2966 ( .A1(byp_alu_rs1_data_e[59]), .A2(n2745), .B(n2678), .Z(
        n3380) );
  HDAOI211D2 U2967 ( .A1(ecl_shft_shift4_e[0]), .A2(n2508), .B(n2302), .C(
        n2303), .Z(n2206) );
  HDEXOR2D1 U2968 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[43]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_11_) );
  HDINVD4 U2969 ( .A(n1773), .Z(n2682) );
  HDNOR3D2 U2970 ( .A1(n2603), .A2(n2604), .A3(n2605), .Z(n2602) );
  HDEXOR2D1 U2971 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[36]), .Z(
        n2127) );
  HDOA21M20D2 U2972 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n91), 
        .A2(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n3), .B(n2128), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n90) );
  HDOA21D1 U2973 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n162), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n93), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n94), .Z(n2128) );
  HDNOR2M1D2 U2974 ( .A1(n3364), .A2(n2200), .Z(n3138) );
  HDOA211D2 U2975 ( .A1(n2912), .A2(n2704), .B(n2853), .C(n2852), .Z(n2893) );
  HDOA211D2 U2976 ( .A1(n2912), .A2(n2456), .B(n2911), .C(n2910), .Z(n2965) );
  HDOA211D2 U2977 ( .A1(n3158), .A2(n2707), .B(n3047), .C(n3046), .Z(n3093) );
  HDOR3DL U2978 ( .A1(n3025), .A2(ecl_alu_out_sel_shift_e_l), .A3(n3576), .Z(
        n2563) );
  HDOR2DL U2979 ( .A1(n2893), .A2(n3576), .Z(n2542) );
  HDAO21D1 U2980 ( .A1(n2481), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n125), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n126), .Z(n2129) );
  HDINVD2 U2981 ( .A(n2695), .Z(n2694) );
  HDEXOR2D1 U2982 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[24]), .Z(
        n2131) );
  HDEXOR2D1 U2983 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[24]), .Z(
        n2130) );
  HDEXOR2D1 U2984 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[24]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I2_24_) );
  HDOAI21DL U2985 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n739), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n712), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n713), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n711) );
  HDNOR3D2 U2986 ( .A1(n2523), .A2(n2524), .A3(n2525), .Z(n2515) );
  HDNOR2M1D2 U2987 ( .A1(n2132), .A2(n2242), .Z(n2239) );
  HDAOI21DL U2988 ( .A1(n2127), .A2(n2240), .B(n2241), .Z(n2132) );
  HDNOR2D2 U2989 ( .A1(n2124), .A2(n2704), .Z(n2208) );
  HDOA21D1 U2990 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n332), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n301), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n302), .Z(n2133) );
  HDEXOR2D1 U2991 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n290), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n20), .Z(alu_adder_out[48])
         );
  HDINVDL U2992 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n668), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n982) );
  HDINVBD4 U2993 ( .A(n2695), .Z(n2299) );
  HDOAI211D2 U2994 ( .A1(n3239), .A2(n2200), .B(n3260), .C(n3238), .Z(n3373)
         );
  HDOAI22M10D1 U2995 ( .A1(ecl_shft_shift4_e[1]), .A2(n2205), .B1(n2300), .B2(
        n2456), .Z(n2329) );
  HDEXNOR2D1 U2996 ( .A1(n1873), .A2(byp_alu_rs2_data_e[32]), .Z(n2136) );
  HDNOR2D4 U2997 ( .A1(n2199), .A2(n2198), .Z(n2138) );
  HDINVD1 U2998 ( .A(n1779), .Z(n2139) );
  HDNOR2D2 U2999 ( .A1(n2663), .A2(n2140), .Z(n2759) );
  HDNOR2M1D1 U3000 ( .A1(n2217), .A2(n2213), .Z(n2210) );
  HDEXOR2D1 U3001 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[35]), .Z(
        n2141) );
  HDNAN3D2 U3002 ( .A1(n2190), .A2(n2431), .A3(n1771), .Z(n2415) );
  HDOAI211D2 U3003 ( .A1(n3198), .A2(n1773), .B(n3260), .C(n3197), .Z(n3354)
         );
  HDAO21DL U3004 ( .A1(n2494), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n491), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n474), .Z(n2142) );
  HDINVD2 U3005 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n476), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n474) );
  HDNAN2D1 U3006 ( .A1(n2395), .A2(n2314), .Z(n2312) );
  HDINVD1 U3007 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n260), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n258) );
  HDAOI21D2 U3008 ( .A1(n2681), .A2(n3283), .B(n3009), .Z(n3200) );
  HDAOI22M20D1 U3009 ( .B1(n2612), .B2(n1924), .A1(n2689), .A2(n2144), .Z(
        n2606) );
  HDOR2D2 U3010 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_17_), .A2(
        byp_alu_rs1_data_e[49]), .Z(n2485) );
  HDAOI22DL U3011 ( .A1(ecl_shft_shift4_e[2]), .A2(n3570), .B1(n2502), .B2(
        ecl_shft_shift4_e[1]), .Z(n2263) );
  HDEXOR2D1 U3012 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[15]), .Z(
        n2146) );
  HDEXOR2D1 U3013 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[18]), .Z(
        n2147) );
  HDOAI22D1 U3014 ( .A1(n2149), .A2(n2689), .B1(n2214), .B2(
        ecl_alu_out_sel_shift_e_l), .Z(n2213) );
  HDNAN2D2 U3015 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n715), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n692), .Z(n2498) );
  HDOR2D2 U3016 ( .A1(n1743), .A2(n2152), .Z(n3362) );
  HDOA21M20D2 U3017 ( .A1(n2486), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n423), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n408), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n404) );
  HDNAN2D2 U3018 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_22_), 
        .A2(byp_alu_rs1_data_e[54]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n175) );
  HDINVD2 U3019 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n430), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n432) );
  HDOR2D4 U3020 ( .A1(n1743), .A2(n2154), .Z(n3381) );
  HDOAI21DL U3021 ( .A1(n1868), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n778), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n773), .Z(n2155) );
  HDNAN2D2 U3022 ( .A1(n2171), .A2(byp_alu_rs1_data_e[20]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n773) );
  HDOAI21M20D2 U3023 ( .A1(n1782), .A2(n3418), .B(n2657), .Z(n3528) );
  HDOA211D4 U3024 ( .A1(n3383), .A2(n2685), .B(n2734), .C(n3381), .Z(n2887) );
  HDINVBD4 U3025 ( .A(n1776), .Z(n2684) );
  HDINVD4 U3026 ( .A(n3528), .Z(n3454) );
  HDAOI21D4 U3027 ( .A1(n1782), .A2(n3380), .B(n3379), .Z(n3493) );
  HDOAI22DL U3028 ( .A1(n3270), .A2(n2702), .B1(n3269), .B2(n3533), .Z(n3273)
         );
  HDOAI22DL U3029 ( .A1(n3270), .A2(n3560), .B1(n3269), .B2(n3563), .Z(n3229)
         );
  HDOAI22DL U3030 ( .A1(n3270), .A2(n3561), .B1(n3269), .B2(n1789), .Z(n3208)
         );
  HDOAI22M10D1 U3031 ( .A1(ecl_shft_shift4_e[0]), .A2(n3514), .B1(n2704), .B2(
        n3478), .Z(n3404) );
  HDEXOR2D1 U3032 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[34]), .Z(
        n2157) );
  HDAOI22DL U3033 ( .A1(n2116), .A2(n3152), .B1(n3151), .B2(
        byp_alu_rs1_data_e[26]), .Z(n3154) );
  HDINVDL U3034 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n694), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n984) );
  HDOAI21DL U3035 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n739), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n660), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n661), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n659) );
  HDAOI21DL U3036 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n689), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n983), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n676), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n674) );
  HDEXOR2D1 U3037 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[5]), .Z(
        n2159) );
  HDEXOR2D1 U3038 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[21]), .Z(
        n2161) );
  HDEXOR2D1 U3039 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[21]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I2_21_) );
  HDNOR2D4 U3040 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n89), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n72), .Z(n2292) );
  HDNAN2D2 U3041 ( .A1(ifu_exu_invert_d), .A2(n2164), .Z(n2165) );
  HDNAN2D2 U3042 ( .A1(n2165), .A2(n2166), .Z(alu_addsub_rs2_data[13]) );
  HDOAI21DL U3043 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n739), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n725), .B(n2134), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n724) );
  HDNAN2D1 U3044 ( .A1(alu_addsub_rs2_data[13]), .A2(byp_alu_rs1_data_e[13]), 
        .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n855) );
  HDAOI31M10D1 U3045 ( .A1(n2283), .A2(n2281), .A3(n2279), .B(n2282), .Z(n2277) );
  HDNOR3D2 U3046 ( .A1(n2582), .A2(n2581), .A3(n1972), .Z(n2580) );
  HDINVBD4 U3047 ( .A(n2679), .Z(n2678) );
  HDEXOR2D1 U3048 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[12]), .Z(
        n2168) );
  HDAOI22DL U3049 ( .A1(n2695), .A2(n3237), .B1(n3536), .B2(n3407), .Z(n2713)
         );
  HDAOI22D1 U3050 ( .A1(n1786), .A2(n3080), .B1(n3536), .B2(n3318), .Z(n2733)
         );
  HDEXOR2D1 U3051 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[20]), .Z(
        n2171) );
  HDAOI21D1 U3052 ( .A1(n2697), .A2(n3258), .B(n3413), .Z(n2729) );
  HDEXOR2D1 U3053 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[11]), .Z(
        n2173) );
  HDEXOR2D1 U3054 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[14]), .Z(
        n2174) );
  HDEXOR2D1 U3055 ( .A1(byp_alu_rs2_data_e[4]), .A2(ifu_exu_invert_d), .Z(
        n2331) );
  HDOA211D2 U3056 ( .A1(n3316), .A2(n2299), .B(n2236), .C(n3315), .Z(n3421) );
  HDOA211D2 U3057 ( .A1(n3566), .A2(n3422), .B(n2367), .C(n2368), .Z(n2369) );
  HDINVD2 U3058 ( .A(n1768), .Z(n2662) );
  HDEXOR2D1 U3059 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[22]), .Z(
        n2179) );
  HDINVD2 U3060 ( .A(n3001), .Z(n2180) );
  HDNOR4D1 U3061 ( .A1(n2184), .A2(n3189), .A3(n3188), .A4(n3187), .Z(n3195)
         );
  HDOAI22D1 U3062 ( .A1(n2924), .A2(n1783), .B1(n2923), .B2(n3576), .Z(n2915)
         );
  HDINVD1 U3063 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n989), .Z(
        n2185) );
  HDINVD2 U3064 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n412), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n587) );
  HDNOR2D2 U3065 ( .A1(n2654), .A2(n3422), .Z(n3266) );
  HDEXOR2D1 U3066 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[41]), .Z(
        n2187) );
  HDNOR2D2 U3067 ( .A1(n3110), .A2(n3109), .Z(n3157) );
  HDNAN2D2 U3068 ( .A1(n2743), .A2(byp_alu_rs1_data_e[8]), .Z(n3498) );
  HDOAI22M10D1 U3069 ( .A1(ecl_shft_shift4_e[0]), .A2(n3302), .B1(n3335), .B2(
        n2704), .Z(n2307) );
  HDNAN2DL U3070 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n989), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n752), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n606) );
  HDNOR2D2 U3071 ( .A1(n2360), .A2(ecl_shft_op32_e), .Z(n2198) );
  HDOAI22D1 U3072 ( .A1(n3205), .A2(n3561), .B1(n3204), .B2(n1789), .Z(n3146)
         );
  HDOAI22M10DL U3073 ( .A1(n1787), .A2(n3204), .B1(n3205), .B2(n2702), .Z(
        n3206) );
  HDNOR4M1D1 U3074 ( .A1(n2188), .A2(n3168), .A3(n3167), .A4(n3166), .Z(n3174)
         );
  HDOA22D1 U3075 ( .A1(n3157), .A2(n3533), .B1(n3156), .B2(n2702), .Z(n2188)
         );
  HDINVD1 U3076 ( .A(n2675), .Z(n2304) );
  HDOAI21D1 U3077 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n366), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n331), .B(n2191), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n330) );
  HDAOI21D4 U3078 ( .A1(n2680), .A2(n3370), .B(n3160), .Z(n3335) );
  HDAOI22D1 U3079 ( .A1(n1786), .A2(n3318), .B1(n2680), .B2(n3080), .Z(n2819)
         );
  HDAOI21DL U3080 ( .A1(n2493), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n355), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n338), .Z(n2191) );
  HDNAN2D1 U3081 ( .A1(n2163), .A2(n2393), .Z(n2376) );
  HDINVDL U3082 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n854), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n997) );
  HDINVDL U3083 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n403), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n397) );
  HDOAI21M20D2 U3084 ( .A1(byp_alu_rs1_data_e[57]), .A2(n2745), .B(n2659), .Z(
        n3364) );
  HDOAI21M20D1 U3085 ( .A1(byp_alu_rs1_data_e[36]), .A2(n2745), .B(n2659), .Z(
        n3080) );
  HDEXOR2D1 U3086 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[42]), .Z(
        alu_addsub_rs2_data[42]) );
  HDINVDL U3087 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n847), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n996) );
  HDINVDL U3088 ( .A(n2332), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n866) );
  HDINVDL U3089 ( .A(n2469), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n561) );
  HDAOI22DL U3090 ( .A1(n2159), .A2(n2828), .B1(n2827), .B2(
        byp_alu_rs1_data_e[5]), .Z(n2830) );
  HDAOI211D4 U3091 ( .A1(ecl_shft_shift4_e[1]), .A2(n3373), .B(n3338), .C(
        n3337), .Z(n3369) );
  HDNAN2D2 U3092 ( .A1(n1742), .A2(n2201), .Z(n2361) );
  HDNOR2D2 U3093 ( .A1(ecl_shft_op32_e), .A2(byp_alu_rs2_data_e[4]), .Z(n2201)
         );
  HDOAI211D1 U3094 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n158), 
        .A2(n2340), .B(n2344), .C(n2345), .Z(n2355) );
  HDAOI21D2 U3095 ( .A1(n2480), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n159), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n160), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n158) );
  HDNAN2D1 U3096 ( .A1(n2163), .A2(n2292), .Z(n2279) );
  HDNAN2DL U3097 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n997), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n855), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n614) );
  HDINVD4 U3098 ( .A(n2202), .Z(n2701) );
  HDAOI22D1 U3099 ( .A1(n3536), .A2(n3535), .B1(n2698), .B2(
        byp_alu_rs1_data_e[61]), .Z(n3537) );
  HDNAN2M1D1 U3100 ( .A1(n3355), .A2(n2699), .Z(n3357) );
  HDNAN2M1D1 U3101 ( .A1(n3346), .A2(n2203), .Z(n3348) );
  HDAND2D1 U3102 ( .A1(n2138), .A2(byp_alu_rs1_data_e[27]), .Z(n3163) );
  HDAOI22D1 U3103 ( .A1(n3536), .A2(n3474), .B1(n2701), .B2(
        byp_alu_rs1_data_e[54]), .Z(n3475) );
  HDAOI22D1 U3104 ( .A1(n3536), .A2(n3483), .B1(n2700), .B2(
        byp_alu_rs1_data_e[55]), .Z(n3484) );
  HDAOI22D1 U3105 ( .A1(n3536), .A2(n3464), .B1(n2700), .B2(
        byp_alu_rs1_data_e[53]), .Z(n3465) );
  HDAOI21M20D2 U3106 ( .A1(n3553), .A2(n1773), .B(n2204), .Z(n2205) );
  HDOAI22D1 U3107 ( .A1(n3332), .A2(n2710), .B1(n2205), .B2(n2705), .Z(n2303)
         );
  HDOAI22D1 U3108 ( .A1(n3334), .A2(n2702), .B1(n2206), .B2(n3563), .Z(n2428)
         );
  HDNOR2D2 U3109 ( .A1(n2360), .A2(ecl_shft_op32_e), .Z(n2207) );
  HDMUXB2DL U3110 ( .A0(n1772), .A1(n1767), .SL(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_17_), .Z(n2215) );
  HDINVD1 U3111 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n4), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n293) );
  HDAOI21D1 U3112 ( .A1(n2215), .A2(n1769), .B(n2216), .Z(n2212) );
  HDOAI21D1 U3113 ( .A1(n2703), .A2(byp_alu_rs1_data_e[49]), .B(n1769), .Z(
        n2211) );
  HDAOI21DL U3114 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_17_), 
        .A2(n2211), .B(n2212), .Z(n2217) );
  HDAOI21D1 U3115 ( .A1(n2013), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n274), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n275), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n273) );
  HDOAI21M20D1 U3116 ( .A1(alu_adder_out_49_), .A2(n1785), .B(n2210), .Z(
        alu_byp_rd_data_e[49]) );
  HDOAI211D1 U3117 ( .A1(n2218), .A2(n2219), .B(n2220), .C(n2221), .Z(
        alu_byp_rd_data_e[54]) );
  HDNAN2M1D1 U3118 ( .A1(n2689), .A2(byp_alu_rs2_data_e[54]), .Z(n2224) );
  HDOAI21D1 U3119 ( .A1(n2703), .A2(byp_alu_rs1_data_e[54]), .B(n1769), .Z(
        n2225) );
  HDNOR4D1 U3120 ( .A1(n2228), .A2(n2229), .A3(n2230), .A4(n2231), .Z(n2222)
         );
  HDOAI22D1 U3121 ( .A1(n3491), .A2(n3576), .B1(n3490), .B2(n1783), .Z(n2231)
         );
  HDOAI22D1 U3122 ( .A1(n3501), .A2(n3561), .B1(n3500), .B2(n1789), .Z(n2230)
         );
  HDOAI22D1 U3123 ( .A1(n3492), .A2(n3560), .B1(n2591), .B2(n3563), .Z(n2229)
         );
  HDOAI22D1 U3124 ( .A1(n3471), .A2(n2702), .B1(n3470), .B2(n3533), .Z(n2228)
         );
  HDNAN4D1 U3125 ( .A1(n2218), .A2(n1785), .A3(n2232), .A4(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n192), .Z(n2220) );
  HDOA211D1 U3126 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n192), .A2(
        n2219), .B(n2223), .C(n2224), .Z(n2234) );
  HDNOR2D2 U3127 ( .A1(n2235), .A2(ecl_shft_enshift_e_l), .Z(n3458) );
  HDNAN2D1 U3128 ( .A1(n2699), .A2(byp_alu_rs1_data_e[36]), .Z(n2236) );
  HDOAI22D1 U3129 ( .A1(n3421), .A2(n2456), .B1(n2661), .B2(n2704), .Z(n2238)
         );
  HDNOR2D1 U3130 ( .A1(n3349), .A2(n2706), .Z(n2237) );
  HDOAI22D1 U3131 ( .A1(n3324), .A2(n3576), .B1(n2301), .B2(n1783), .Z(n2245)
         );
  HDOAI22D1 U3132 ( .A1(n3326), .A2(n3560), .B1(n3325), .B2(n3563), .Z(n2246)
         );
  HDOAI22D1 U3133 ( .A1(n3310), .A2(n2702), .B1(n3309), .B2(n3533), .Z(n2244)
         );
  HDNOR3M1D2 U3134 ( .A1(n2249), .A2(n2244), .A3(n1777), .Z(n2243) );
  HDAOI21D1 U3135 ( .A1(n2247), .A2(n1769), .B(n2248), .Z(n2241) );
  HDOAI21D1 U3136 ( .A1(n2703), .A2(byp_alu_rs1_data_e[36]), .B(n1769), .Z(
        n2240) );
  HDOAI21M20D1 U3137 ( .A1(alu_adder_out_36_), .A2(n1785), .B(n2239), .Z(
        alu_byp_rd_data_e[36]) );
  HDNAN4D1 U3138 ( .A1(n2250), .A2(n2251), .A3(n2252), .A4(n2253), .Z(
        alu_byp_rd_data_e[63]) );
  HDAOI21D1 U3139 ( .A1(n2254), .A2(n2255), .B(n2256), .Z(n2253) );
  HDOAI31D1 U3140 ( .A1(n2258), .A2(n2259), .A3(n2260), .B(n2261), .Z(n2252)
         );
  HDAOI21D1 U3141 ( .A1(n2262), .A2(ecl_shft_lshift_e_l), .B(
        ecl_alu_out_sel_shift_e_l), .Z(n2261) );
  HDOAI21M10D1 U3142 ( .A1(ecl_shft_shift1_e[2]), .A2(n3572), .B(n2262), .Z(
        n2260) );
  HDNAN4D1 U3143 ( .A1(n2265), .A2(n1785), .A3(n2266), .A4(n2267), .Z(n2251)
         );
  HDINVBD2 U3144 ( .A(n2254), .Z(n2267) );
  HDAOI211D1 U3145 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n96), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n48), .B(n2269), .C(n2270), 
        .Z(n2268) );
  HDOAI21D1 U3146 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n56), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n50), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n51), .Z(n2269) );
  HDOR2D1 U3147 ( .A1(n2265), .A2(n2271), .Z(n2250) );
  HDNAN3D1 U3148 ( .A1(n2163), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n44), .A3(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n4), .Z(n2265) );
  HDNOR2D2 U3149 ( .A1(n1996), .A2(byp_alu_rs1_data_e[1]), .Z(n2272) );
  HDINVDL U3150 ( .A(n2272), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n1009) );
  HDAOI22D1 U3151 ( .A1(n2274), .A2(n2900), .B1(n2899), .B2(
        byp_alu_rs1_data_e[10]), .Z(n2902) );
  HDNOR2D2 U3152 ( .A1(n2273), .A2(byp_alu_rs1_data_e[10]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n891) );
  HDEXOR2D1 U3153 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[10]), .Z(
        n2273) );
  HDNOR2D2 U3154 ( .A1(alu_addsub_rs2_data[16]), .A2(byp_alu_rs1_data_e[16]), 
        .Z(n2275) );
  HDINVDL U3155 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n891), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n1000) );
  HDNAN2D2 U3156 ( .A1(n2309), .A2(n1865), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n883) );
  HDOAI211D1 U3157 ( .A1(n2276), .A2(ecl_alu_out_sel_shift_e_l), .B(n2278), 
        .C(n2277), .Z(alu_byp_rd_data_e[61]) );
  HDAOI31D1 U3158 ( .A1(n2287), .A2(n2288), .A3(n1769), .B(n2289), .Z(n2286)
         );
  HDNAN2M1D1 U3159 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_29_), 
        .A2(n1772), .Z(n2287) );
  HDNOR2M1D1 U3160 ( .A1(byp_alu_rs2_data_e[61]), .A2(n2689), .Z(n2285) );
  HDOAI21D1 U3161 ( .A1(byp_alu_rs1_data_e[61]), .A2(n2703), .B(n1769), .Z(
        n2284) );
  HDOAI21D1 U3162 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n90), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n72), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n73), .Z(n2283) );
  HDNOR4D1 U3163 ( .A1(n2293), .A2(n2294), .A3(n2295), .A4(n2296), .Z(n2276)
         );
  HDOAI22D1 U3164 ( .A1(n3572), .A2(n1789), .B1(n3573), .B2(n3563), .Z(n2295)
         );
  HDOAI22D1 U3165 ( .A1(n3575), .A2(n3561), .B1(n3534), .B2(n3533), .Z(n2294)
         );
  HDOAI22D1 U3166 ( .A1(n3574), .A2(n3560), .B1(n3544), .B2(n1783), .Z(n2293)
         );
  HDAO21M10D1 U3167 ( .A2(n2283), .A1(n2280), .B(n2297), .Z(n2282) );
  HDNAN2D2 U3168 ( .A1(n2682), .A2(n3143), .Z(n2298) );
  HDNOR2M1D1 U3169 ( .A1(n2695), .A2(n2788), .Z(n2714) );
  HDOA211D4 U3170 ( .A1(n3261), .A2(n2299), .B(n3242), .C(n3002), .Z(n3179) );
  HDOA21M20D2 U3171 ( .A1(n2138), .A2(byp_alu_rs1_data_e[34]), .B(n2362), .Z(
        n2300) );
  HDNOR2D1 U3172 ( .A1(n2300), .A2(n2704), .Z(n2302) );
  HDNOR2D1 U3173 ( .A1(n2300), .A2(n2710), .Z(n3405) );
  HDOA21M20D2 U3174 ( .A1(n1782), .A2(n3100), .B(n2305), .Z(n3302) );
  HDNOR2D1 U3175 ( .A1(n3408), .A2(n2710), .Z(n2306) );
  HDNOR2D2 U3176 ( .A1(n2159), .A2(byp_alu_rs1_data_e[5]), .Z(n2308) );
  HDNOR2D2 U3177 ( .A1(n1781), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n916), .Z(n2309) );
  HDOR2DL U3178 ( .A1(n1781), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n916), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n905) );
  HDNOR2M1D1 U3179 ( .A1(n1792), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n191), .Z(n2314) );
  HDAO21D1 U3180 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n793), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n766), .B(n2155), .Z(n2315)
         );
  HDMUXB2DL U3181 ( .A0(n1772), .A1(n1767), .SL(n1804), .Z(n2322) );
  HDNAN2D1 U3182 ( .A1(n2322), .A2(n1769), .Z(n2321) );
  HDOAI21D1 U3183 ( .A1(n2703), .A2(byp_alu_rs1_data_e[22]), .B(n1769), .Z(
        n2320) );
  HDOAI22D1 U3184 ( .A1(n3104), .A2(n1783), .B1(n3103), .B2(n3576), .Z(n2326)
         );
  HDOAI22D1 U3185 ( .A1(n3094), .A2(n3533), .B1(n3093), .B2(n2702), .Z(n2325)
         );
  HDOAI22D1 U3186 ( .A1(n3118), .A2(n1789), .B1(n3117), .B2(n3561), .Z(n2324)
         );
  HDOAI22D1 U3187 ( .A1(n3106), .A2(n3563), .B1(n3105), .B2(n3560), .Z(n2323)
         );
  HDAOI22D1 U3188 ( .A1(byp_alu_rs2_data_e[22]), .A2(n2683), .B1(
        alu_adder_out_22_), .B2(n1785), .Z(n2319) );
  HDAOI22D1 U3189 ( .A1(n2178), .A2(n2320), .B1(n2321), .B2(
        byp_alu_rs1_data_e[22]), .Z(n2318) );
  HDNOR4D1 U3190 ( .A1(n2323), .A2(n2324), .A3(n2325), .A4(n2326), .Z(n2317)
         );
  HDOAI21M20DL U3191 ( .A1(n3044), .A2(n2684), .B(n3260), .Z(n2327) );
  HDAOI22D1 U3192 ( .A1(n2813), .A2(n2000), .B1(n2812), .B2(
        byp_alu_rs1_data_e[4]), .Z(n2815) );
  HDNAN2D2 U3193 ( .A1(n2331), .A2(byp_alu_rs1_data_e[4]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n951) );
  HDNOR2D2 U3194 ( .A1(n2330), .A2(byp_alu_rs1_data_e[4]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n950) );
  HDOAI21D1 U3195 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n869), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n881), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n870), .Z(n2332) );
  HDEXOR2D1 U3196 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[12]), .Z(
        alu_addsub_rs2_data[12]) );
  HDAOI22D1 U3197 ( .A1(n2334), .A2(n2798), .B1(n2797), .B2(
        byp_alu_rs1_data_e[3]), .Z(n2800) );
  HDNOR2D2 U3198 ( .A1(n2335), .A2(byp_alu_rs1_data_e[3]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n959) );
  HDEXOR2D1 U3199 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[3]), .Z(
        n2333) );
  HDEXOR2D1 U3200 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[3]), .Z(
        n2335) );
  HDOAI21DL U3201 ( .A1(n2464), .A2(n1810), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n951), .Z(n2477) );
  HDINVD1 U3202 ( .A(n1810), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n954) );
  HDNAN2M1D1 U3203 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n447), 
        .A2(n2492), .Z(n2337) );
  HDOAI21D1 U3204 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n532), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n505), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n506), .Z(n2336) );
  HDOAI21D1 U3205 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n430), .A2(
        n2005), .B(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n298), .Z(n2480)
         );
  HDNAN2D1 U3206 ( .A1(n2701), .A2(byp_alu_rs1_data_e[45]), .Z(n2339) );
  HDOAI211D1 U3207 ( .A1(n2341), .A2(n2340), .B(n2342), .C(n2343), .Z(
        alu_byp_rd_data_e[56]) );
  HDNAN2M1D1 U3208 ( .A1(n2689), .A2(byp_alu_rs2_data_e[56]), .Z(n2345) );
  HDAOI22D1 U3209 ( .A1(byp_alu_rs1_data_e[56]), .A2(n2346), .B1(n2347), .B2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_24_), .Z(n2344) );
  HDOAI21D1 U3210 ( .A1(n2703), .A2(byp_alu_rs1_data_e[56]), .B(n1769), .Z(
        n2347) );
  HDOAI211D1 U3211 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_24_), 
        .A2(n2703), .B(n2348), .C(n1769), .Z(n2346) );
  HDOAI31D1 U3212 ( .A1(n2350), .A2(n2351), .A3(n2352), .B(n1924), .Z(n2342)
         );
  HDOAI22D1 U3213 ( .A1(n3501), .A2(n3576), .B1(n3492), .B2(n2702), .Z(n2354)
         );
  HDNAN2M1D1 U3214 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n157), 
        .A2(n2163), .Z(n2341) );
  HDAOI21M10D1 U3215 ( .A1(n2356), .A2(n2341), .B(n2355), .Z(n2343) );
  HDNOR2D2 U3216 ( .A1(n2358), .A2(n2364), .Z(n2359) );
  HDNOR2D2 U3217 ( .A1(n2158), .A2(ecl_shft_op32_e), .Z(n2660) );
  HDINVBD20 U3218 ( .A(n2361), .Z(n2695) );
  HDOAI211D1 U3219 ( .A1(n2365), .A2(n2433), .B(n2434), .C(n2366), .Z(
        alu_byp_rd_data_e[33]) );
  HDAO21M20D1 U3220 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n926), 
        .A2(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n883), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n886), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n882) );
  HDNAN2D2 U3221 ( .A1(alu_addsub_rs2_data[7]), .A2(byp_alu_rs1_data_e[7]), 
        .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n917) );
  HDNAN2D2 U3222 ( .A1(n3550), .A2(byp_alu_rs1_data_e[16]), .Z(n2367) );
  HDOAI22D1 U3223 ( .A1(n2123), .A2(n2710), .B1(n3530), .B2(n2707), .Z(n2371)
         );
  HDNOR2D1 U3224 ( .A1(n3531), .A2(n2704), .Z(n2370) );
  HDAOI21D1 U3225 ( .A1(n1889), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n138), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n139), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n137) );
  HDOAI21M20D1 U3226 ( .A1(alu_adder_out_57_), .A2(n1785), .B(n2372), .Z(
        alu_byp_rd_data_e[57]) );
  HDNOR2D2 U3227 ( .A1(n2173), .A2(byp_alu_rs1_data_e[11]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n880) );
  HDNAN2D2 U3228 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n863), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n845), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n843) );
  HDINVDL U3229 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n883), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n885) );
  HDOAI211D1 U3230 ( .A1(n2376), .A2(n2377), .B(n2378), .C(n2379), .Z(
        alu_byp_rd_data_e[47]) );
  HDAOI211D1 U3231 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_15_), 
        .A2(n2385), .B(n2386), .C(n2387), .Z(n2381) );
  HDNOR2M1D1 U3232 ( .A1(byp_alu_rs2_data_e[47]), .A2(n2689), .Z(n2386) );
  HDOAI21D1 U3233 ( .A1(n2703), .A2(byp_alu_rs1_data_e[47]), .B(n1769), .Z(
        n2385) );
  HDNOR4D1 U3234 ( .A1(n2388), .A2(n2389), .A3(n2390), .A4(n2391), .Z(n2380)
         );
  HDOAI22D1 U3235 ( .A1(n3428), .A2(n3560), .B1(n3427), .B2(n3563), .Z(n2391)
         );
  HDOAI22D1 U3236 ( .A1(n3433), .A2(n3561), .B1(n1994), .B2(n1789), .Z(n2390)
         );
  HDOAI22D1 U3237 ( .A1(n3415), .A2(n3576), .B1(n2590), .B2(n1783), .Z(n2389)
         );
  HDOAI22D1 U3238 ( .A1(n3406), .A2(n2702), .B1(n1779), .B2(n3533), .Z(n2388)
         );
  HDOA21D1 U3239 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n328), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n310), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n311), .Z(n2384) );
  HDNOR2M1D1 U3240 ( .A1(n1791), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n327), .Z(n2393) );
  HDAOI22D1 U3241 ( .A1(n2394), .A2(n2781), .B1(n2780), .B2(
        byp_alu_rs1_data_e[2]), .Z(n2782) );
  HDOAI211D1 U3242 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n362), 
        .A2(n2397), .B(n2401), .C(n2402), .Z(n2400) );
  HDNAN2M1D1 U3243 ( .A1(n2689), .A2(byp_alu_rs2_data_e[44]), .Z(n2402) );
  HDOAI21D1 U3244 ( .A1(byp_alu_rs1_data_e[44]), .A2(n2703), .B(n1769), .Z(
        n2404) );
  HDAOI21D1 U3245 ( .A1(n2407), .A2(n2408), .B(ecl_alu_out_sel_shift_e_l), .Z(
        n2399) );
  HDAOI21M20D1 U3246 ( .A1(n3387), .A2(n3533), .B(n2409), .Z(n2408) );
  HDOAI222D1 U3247 ( .A1(n3406), .A2(n3561), .B1(n3388), .B2(n2702), .C1(n2114), .C2(n3563), .Z(n2409) );
  HDAOI211D1 U3248 ( .A1(n2139), .A2(n2688), .B(n2410), .C(n2411), .Z(n2407)
         );
  HDOAI22D1 U3249 ( .A1(n3395), .A2(n3576), .B1(n3397), .B2(n3560), .Z(n2410)
         );
  HDOAI211D1 U3250 ( .A1(n2414), .A2(n2415), .B(n2417), .C(n2416), .Z(
        alu_byp_rd_data_e[39]) );
  HDAOI211D1 U3251 ( .A1(n2421), .A2(n2182), .B(n2422), .C(n2423), .Z(n2420)
         );
  HDNOR2M1D1 U3252 ( .A1(byp_alu_rs2_data_e[39]), .A2(n2689), .Z(n2423) );
  HDAOI31D1 U3253 ( .A1(n2424), .A2(n1769), .A3(n2425), .B(n3486), .Z(n2422)
         );
  HDNAN2M1D1 U3254 ( .A1(n2182), .A2(n1772), .Z(n2424) );
  HDOAI21D1 U3255 ( .A1(n2703), .A2(byp_alu_rs1_data_e[39]), .B(n1769), .Z(
        n2421) );
  HDNOR4D1 U3256 ( .A1(n2426), .A2(n2427), .A3(n2428), .A4(n2429), .Z(n2418)
         );
  HDOAI22D1 U3257 ( .A1(n3369), .A2(n3561), .B1(n3368), .B2(n1789), .Z(n2429)
         );
  HDNOR2M1D1 U3258 ( .A1(n3562), .A2(n3342), .Z(n2427) );
  HDOAI222D1 U3259 ( .A1(n3361), .A2(n3560), .B1(n3343), .B2(n3576), .C1(n3333), .C2(n3533), .Z(n2426) );
  HDOAI21M20D1 U3260 ( .A1(n2437), .A2(ecl_alu_out_sel_shift_e_l), .B(n2438), 
        .Z(n2434) );
  HDOAI22D1 U3261 ( .A1(n3310), .A2(n3561), .B1(n3309), .B2(n1789), .Z(n2441)
         );
  HDOAI22D1 U3262 ( .A1(n3293), .A2(n1783), .B1(n3294), .B2(n3576), .Z(n2440)
         );
  HDNAN2M1D1 U3263 ( .A1(n2689), .A2(byp_alu_rs2_data_e[33]), .Z(n2444) );
  HDAOI22D1 U3264 ( .A1(byp_alu_rs1_data_e[33]), .A2(n2445), .B1(n2446), .B2(
        n2151), .Z(n2442) );
  HDOAI21D1 U3265 ( .A1(n2703), .A2(byp_alu_rs1_data_e[33]), .B(n1769), .Z(
        n2446) );
  HDNOR2D1 U3266 ( .A1(n2440), .A2(n2441), .Z(n2439) );
  HDEXOR2D1 U3267 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[40]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_8_) );
  HDNAN2D2 U3268 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_8_), .A2(
        byp_alu_rs1_data_e[40]), .Z(n2447) );
  HDNAN2DL U3269 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n587), .A2(
        n2447), .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n28) );
  HDOA211D2 U3270 ( .A1(n3261), .A2(n2200), .B(n3260), .C(n3259), .Z(n3378) );
  HDOA21M20D2 U3271 ( .A1(n3311), .A2(n1782), .B(n2658), .Z(n3416) );
  HDNAN2DL U3272 ( .A1(ecl_shft_shift4_e[2]), .A2(n3457), .Z(n2450) );
  HDNOR2D2 U3273 ( .A1(n2451), .A2(byp_alu_rs1_data_e[48]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n276) );
  HDNAN2D2 U3274 ( .A1(n1977), .A2(byp_alu_rs1_data_e[48]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n277) );
  HDAO21M20DL U3275 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n739), 
        .A2(n2112), .B(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n689), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n685) );
  HDAOI22M10D1 U3276 ( .B1(alu_adder_out[27]), .B2(n1785), .A1(n2452), .A2(
        n2683), .Z(n3172) );
  HDEXNOR2DL U3277 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n596), 
        .A2(n2479), .Z(alu_adder_out[31]) );
  HDINVDL U3278 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n268), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n262) );
  HDEXOR2D2 U3279 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[51]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_19_) );
  HDAOI211D1 U3280 ( .A1(n3018), .A2(n3445), .B(n2979), .C(n2978), .Z(n2453)
         );
  HDOAI22M10D1 U3281 ( .A1(n3562), .A2(n3026), .B1(n3058), .B2(n1789), .Z(
        n2573) );
  HDOAI22D1 U3282 ( .A1(n2977), .A2(n3565), .B1(n3521), .B2(n3040), .Z(n2978)
         );
  HDOA22D1 U3283 ( .A1(n2837), .A2(n1783), .B1(n2817), .B2(n2702), .Z(n2468)
         );
  HDINVD2 U3284 ( .A(n3165), .Z(n3018) );
  HDNOR2D2 U3285 ( .A1(n2717), .A2(ecl_shft_enshift_e_l), .Z(n3474) );
  HDOAI21M20D2 U3286 ( .A1(n3474), .A2(n2681), .B(n3085), .Z(n3298) );
  HDNAN2DL U3287 ( .A1(n2701), .A2(byp_alu_rs1_data_e[57]), .Z(n3504) );
  HDINVD4 U3288 ( .A(n3096), .Z(n2959) );
  HDOR2D1 U3289 ( .A1(n2360), .A2(ecl_shft_op32_e), .Z(n2454) );
  HDAOI22D1 U3290 ( .A1(n1786), .A2(n3389), .B1(n2682), .B2(n3196), .Z(n2945)
         );
  HDINVBD2 U3291 ( .A(n3547), .Z(n3544) );
  HDAOI211D2 U3292 ( .A1(n3018), .A2(n3474), .B(n3017), .C(n3016), .Z(n3076)
         );
  HDOA211D2 U3293 ( .A1(n3305), .A2(n2694), .B(n3304), .C(n3303), .Z(n3411) );
  HDAOI22M10D1 U3294 ( .B1(ecl_shft_shift4_e[2]), .B2(n3011), .A1(n2710), .A2(
        n3084), .Z(n2885) );
  HDNOR2D2 U3295 ( .A1(n2753), .A2(n2666), .Z(n2755) );
  HDNOR2D2 U3296 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n694), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n707), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n692) );
  HDNOR2D2 U3297 ( .A1(n2006), .A2(byp_alu_rs1_data_e[25]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n707) );
  HDNOR2D2 U3298 ( .A1(n3141), .A2(n3140), .Z(n3205) );
  HDAOI211D2 U3299 ( .A1(ecl_shft_shift4_e[1]), .A2(n3298), .B(n3145), .C(
        n3144), .Z(n3204) );
  HDINVD2 U3300 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n514), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n593) );
  HDINVDL U3301 ( .A(n1814), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n896) );
  HDNAN2D2 U3302 ( .A1(n2161), .A2(byp_alu_rs1_data_e[21]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n752) );
  HDOAI21M20D2 U3303 ( .A1(byp_alu_rs1_data_e[56]), .A2(n2745), .B(n2678), .Z(
        n1756) );
  HDNAN2D2 U3304 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n591), .A2(
        n2494), .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n471) );
  HDOAI22D1 U3305 ( .A1(n3374), .A2(n2456), .B1(n3341), .B2(n2704), .Z(n3243)
         );
  HDOAI21M20D1 U3306 ( .A1(alu_adder_out[60]), .A2(n1785), .B(n2643), .Z(
        alu_byp_rd_data_e[60]) );
  HDNAN3D2 U3307 ( .A1(n2458), .A2(n2543), .A3(n2542), .Z(n2544) );
  HDAOI21D2 U3308 ( .A1(n2682), .A2(n3318), .B(n3081), .Z(n3284) );
  HDINVDL U3309 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n751), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n989) );
  HDNAN3D2 U3310 ( .A1(n2776), .A2(n3005), .A3(n2961), .Z(n2962) );
  HDNOR2D2 U3311 ( .A1(n2671), .A2(ecl_alu_out_sel_shift_e_l), .Z(n2663) );
  HDOAI222D1 U3312 ( .A1(n2807), .A2(n3563), .B1(n3576), .B2(n1733), .C1(n1789), .C2(n2822), .Z(n2779) );
  HDINVD4 U3313 ( .A(n1778), .Z(n2653) );
  HDOA22D2 U3314 ( .A1(n3428), .A2(n3576), .B1(n3427), .B2(n1783), .Z(n2462)
         );
  HDAOI211D2 U3315 ( .A1(ecl_shft_shift4_e[1]), .A2(n3543), .B(n3542), .C(
        n3541), .Z(n3572) );
  HDINVDL U3316 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n959), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n953) );
  HDNAN2D2 U3317 ( .A1(n2127), .A2(byp_alu_rs1_data_e[36]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n481) );
  HDNOR2D2 U3318 ( .A1(n3007), .A2(n3006), .Z(n3058) );
  HDNOR3D4 U3319 ( .A1(n2927), .A2(n3163), .A3(n2181), .Z(n3111) );
  HDAOI21D4 U3320 ( .A1(n1782), .A2(n3370), .B(n3379), .Z(n3481) );
  HDINVD2 U3321 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n481), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n491) );
  HDINVDL U3322 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n364), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n366) );
  HDNAN2D2 U3323 ( .A1(alu_addsub_rs2_data[38]), .A2(byp_alu_rs1_data_e[38]), 
        .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n447) );
  HDEXOR2D2 U3324 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[38]), .Z(
        alu_addsub_rs2_data[38]) );
  HDNOR2D2 U3325 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n127), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n97), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n95) );
  HDOAI21D1 U3326 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n532), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n505), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n506), .Z(n2466) );
  HDNAN2D2 U3327 ( .A1(n1869), .A2(n2490), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n369) );
  HDNAN2D2 U3328 ( .A1(n2690), .A2(byp_alu_rs1_data_e[29]), .Z(n3393) );
  HDINVD4 U3329 ( .A(n1744), .Z(n2690) );
  HDNAN2D2 U3330 ( .A1(n2131), .A2(byp_alu_rs1_data_e[24]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n721) );
  HDOA211D4 U3331 ( .A1(n3394), .A2(n2685), .B(n2742), .C(n3393), .Z(n2892) );
  HDAOI21D1 U3332 ( .A1(n2485), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n287), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n270), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n268) );
  HDAOI211D2 U3333 ( .A1(ecl_shft_shift4_e[1]), .A2(n2775), .B(n2750), .C(
        n2749), .Z(n2766) );
  HDNAN2D2 U3334 ( .A1(n1981), .A2(byp_alu_rs1_data_e[44]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n345) );
  HDOA211D2 U3335 ( .A1(n2887), .A2(n2456), .B(n2886), .C(n2885), .Z(n2923) );
  HDNAN2D2 U3336 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n593), .A2(
        n1770), .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n505) );
  HDNOR4M1D1 U3337 ( .A1(n2468), .A2(n2825), .A3(n2823), .A4(n2824), .Z(n2831)
         );
  HDEXOR2D1 U3338 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[33]), .Z(
        alu_addsub_rs2_data[33]) );
  HDNAN2D2 U3339 ( .A1(n2660), .A2(n3282), .Z(n2470) );
  HDOA21M20D2 U3340 ( .A1(n2478), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n261), .B(n2471), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n260) );
  HDINVDL U3341 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n739), .Z(
        n2472) );
  HDOAI21DL U3342 ( .A1(n2153), .A2(n2134), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n721), .Z(n2473) );
  HDNOR2D2 U3343 ( .A1(alu_addsub_rs2_data[13]), .A2(byp_alu_rs1_data_e[13]), 
        .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n854) );
  HDNAN2D2 U3344 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n577), .A2(
        n2495), .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n233) );
  HDNAN2DL U3345 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n896), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n903), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n618) );
  HDINVD1 U3346 ( .A(n2459), .Z(n2474) );
  HDAOI22DL U3347 ( .A1(n2147), .A2(n3033), .B1(n3032), .B2(
        byp_alu_rs1_data_e[18]), .Z(n3035) );
  HDINVD1 U3348 ( .A(n1793), .Z(n2476) );
  HDAOI211D2 U3349 ( .A1(ecl_shft_shift4_e[2]), .A2(n3510), .B(n3456), .C(
        n3435), .Z(n3469) );
  HDOA211D2 U3350 ( .A1(n3553), .A2(n2694), .B(n3403), .C(n3402), .Z(n3514) );
  HDOAI21D1 U3351 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n720), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n726), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n721), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n715) );
  HDOAI21D1 U3352 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n430), .A2(
        n2005), .B(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n298), .Z(n2478)
         );
  HDOR2D1 U3353 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_15_), .A2(
        byp_alu_rs1_data_e[47]), .Z(n2489) );
  HDOR2D1 U3354 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_19_), .A2(
        byp_alu_rs1_data_e[51]), .Z(n2495) );
  HDOR2D1 U3355 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_21_), .A2(
        byp_alu_rs1_data_e[53]), .Z(n2488) );
  HDINVD1 U3356 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n510), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n508) );
  HDINVD1 U3357 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n311), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n321) );
  HDINVD1 U3358 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n89), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n87) );
  HDOAI21D1 U3359 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n430), .A2(
        n2122), .B(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n298), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n3) );
  HDINVD1 U3360 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n107), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n117) );
  HDINVD1 U3361 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n90), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n88) );
  HDAOI21D1 U3362 ( .A1(n2395), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n87), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n88), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n86) );
  HDINVD1 U3363 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n123), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n121) );
  HDINVD1 U3364 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n471), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n465) );
  HDINVD1 U3365 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n259), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n257) );
  HDAOI21D1 U3366 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n839), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n710), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n711), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n709) );
  HDAOI21D1 U3367 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n839), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n684), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n685), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n683) );
  HDNOR2D2 U3368 ( .A1(alu_addsub_rs2_data[17]), .A2(byp_alu_rs1_data_e[17]), 
        .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n803) );
  HDNOR2D2 U3369 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n777), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n772), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n766) );
  HDNOR2D2 U3370 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I2_21_), 
        .A2(byp_alu_rs1_data_e[21]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n751) );
  HDNAN2D2 U3371 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n766), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n744), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n742) );
  HDNOR2D2 U3372 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I2_24_), 
        .A2(byp_alu_rs1_data_e[24]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n720) );
  HDNOR2D2 U3373 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n725), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n720), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n714) );
  HDNOR2D2 U3374 ( .A1(n2116), .A2(byp_alu_rs1_data_e[26]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n694) );
  HDNAN2D2 U3375 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n714), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n692), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n686) );
  HDNOR2D2 U3376 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I2_29_), 
        .A2(byp_alu_rs1_data_e[29]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n651) );
  HDNOR2D2 U3377 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n638), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n686), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n636) );
  HDNOR2D2 U3378 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_4_), .A2(
        byp_alu_rs1_data_e[36]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n480) );
  HDNAN2D2 U3379 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n499), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n435), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n429) );
  HDNOR2D2 U3380 ( .A1(n1998), .A2(byp_alu_rs1_data_e[9]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n902) );
  HDNOR2D2 U3381 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I2_20_), 
        .A2(byp_alu_rs1_data_e[20]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n772) );
  HDNOR2D2 U3382 ( .A1(n2179), .A2(byp_alu_rs1_data_e[22]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n746) );
  HDNOR2D2 U3383 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n751), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n746), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n744) );
  HDNOR2D2 U3384 ( .A1(n1866), .A2(byp_alu_rs1_data_e[27]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n681) );
  HDNOR2D2 U3385 ( .A1(n1975), .A2(byp_alu_rs1_data_e[28]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n668) );
  HDNOR2D2 U3386 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I2_30_), 
        .A2(byp_alu_rs1_data_e[30]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n642) );
  HDNAN2D2 U3387 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n589), .A2(
        n2492), .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n437) );
  HDNAN2D2 U3388 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n583), .A2(
        n2493), .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n331) );
  HDINVDL U3389 ( .A(n2473), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n713) );
  HDINVD1 U3390 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n687), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n689) );
  HDNOR2D2 U3391 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n798), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n803), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n796) );
  HDINVD1 U3392 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n681), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n983) );
  HDINVD1 U3393 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n880), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n999) );
  HDINVD1 U3394 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n869), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n998) );
  HDINVD1 U3395 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n837), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n995) );
  HDAOI21D1 U3396 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n839), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n736), .B(n2472), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n735) );
  HDINVD1 U3397 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n916), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n1003) );
  HDAOI21D4 U3398 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n228), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n163), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n164), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n162) );
  HDOAI21D1 U3399 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n162), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n127), .B(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n128), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n126) );
  HDNOR2D2 U3400 ( .A1(n2497), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n54), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n52) );
  HDINVD2 U3401 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n446), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n589) );
  HDNOR2D2 U3402 ( .A1(alu_addsub_rs2_data[38]), .A2(byp_alu_rs1_data_e[38]), 
        .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n446) );
  HDNOR2D2 U3403 ( .A1(n2157), .A2(byp_alu_rs1_data_e[34]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n514) );
  HDNOR2D2 U3404 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_22_), 
        .A2(byp_alu_rs1_data_e[54]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n174) );
  HDNAN2D2 U3405 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n575), .A2(
        n2488), .Z(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n195) );
  HDNOR2D2 U3406 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n195), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n165), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n163) );
  HDNAN2D2 U3407 ( .A1(n1792), .A2(n2487), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n165) );
  HDNOR2D2 U3408 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_14_), 
        .A2(byp_alu_rs1_data_e[46]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n310) );
  HDNAN2D2 U3409 ( .A1(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n4), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n91), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n89) );
  HDNAN2D2 U3410 ( .A1(n1791), .A2(n2489), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n301) );
  HDAND2D2 U3411 ( .A1(n2498), .A2(n1780), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_n687) );
  HDINVD2 U3412 ( .A(n1743), .Z(n2691) );
  HDNOR2D2 U3413 ( .A1(n3335), .A2(n2456), .Z(n3338) );
  HDAOI22D1 U3414 ( .A1(n2695), .A2(n3295), .B1(n2680), .B2(n3019), .Z(n2776)
         );
  HDINVBD4 U3415 ( .A(n2695), .Z(n2654) );
  HDOAI21M20D1 U3416 ( .A1(n1782), .A2(n3080), .B(n3260), .Z(n3081) );
  HDAOI21D1 U3417 ( .A1(n1786), .A2(n3301), .B(n3015), .Z(n2787) );
  HDAOI21D2 U3418 ( .A1(n2681), .A2(n3295), .B(n3020), .Z(n3220) );
  HDOAI21M20D1 U3419 ( .A1(n1782), .A2(n3019), .B(n3260), .Z(n3020) );
  HDNAN2DL U3420 ( .A1(n2695), .A2(n3061), .Z(n2723) );
  HDNAN2D1 U3421 ( .A1(n2684), .A2(n3000), .Z(n3242) );
  HDOAI22DL U3422 ( .A1(n2822), .A2(n3563), .B1(n2785), .B2(n2702), .Z(n2796)
         );
  HDNOR2D2 U3423 ( .A1(n2785), .A2(n1795), .Z(n2754) );
  HDNAN2D8 U3424 ( .A1(n2684), .A2(ecl_shft_shift4_e[0]), .Z(n2977) );
  HDNAN2D2 U3425 ( .A1(n2908), .A2(n3445), .Z(n2837) );
  HDNAN2D2 U3426 ( .A1(n2908), .A2(n2888), .Z(n2822) );
  HDINVD4 U3427 ( .A(n3001), .Z(n2961) );
  HDINVD4 U3428 ( .A(n1773), .Z(n2680) );
  HDINVD4 U3429 ( .A(n2744), .Z(n2679) );
  HDOAI21M20D1 U3430 ( .A1(n2684), .A2(n3159), .B(n3260), .Z(n3160) );
  HDNAN2D2 U3431 ( .A1(alu_adder_out[62]), .A2(n1785), .Z(n2607) );
  HDAOI211D2 U3432 ( .A1(byp_alu_rs1_data_e[32]), .A2(n2699), .B(n3266), .C(
        n3265), .Z(n3384) );
  HDAOI21D4 U3433 ( .A1(n1782), .A2(n1756), .B(n3379), .Z(n3462) );
  HDINVD4 U3434 ( .A(n2658), .Z(n3379) );
  HDAOI211D2 U3435 ( .A1(ecl_shft_shift4_e[0]), .A2(n3354), .B(n3353), .C(
        n3352), .Z(n3388) );
  HDOAI21M20D1 U3436 ( .A1(n2684), .A2(n3088), .B(n3260), .Z(n3089) );
  HDOAI21M20D1 U3437 ( .A1(byp_alu_rs1_data_e[37]), .A2(n2745), .B(n2659), .Z(
        n3088) );
  HDOAI22D1 U3438 ( .A1(n2453), .A2(n3563), .B1(n3013), .B2(n1783), .Z(n2556)
         );
  HDAOI22D1 U3439 ( .A1(n2695), .A2(n3112), .B1(n3536), .B2(n3344), .Z(n2730)
         );
  HDAOI22D1 U3440 ( .A1(n3139), .A2(n2695), .B1(n3536), .B2(n3364), .Z(n2746)
         );
  HDNAN2D2 U3441 ( .A1(n2908), .A2(n2866), .Z(n2792) );
  HDAOI22D1 U3442 ( .A1(n2695), .A2(n3159), .B1(n3536), .B2(n3370), .Z(n2719)
         );
  HDAOI22D1 U3443 ( .A1(n1786), .A2(n3100), .B1(n3336), .B2(n3536), .Z(n2718)
         );
  HDAOI22D1 U3444 ( .A1(n2172), .A2(n2919), .B1(n2918), .B2(
        byp_alu_rs1_data_e[11]), .Z(n2921) );
  HDNAN3D1 U3445 ( .A1(n2761), .A2(n2996), .A3(n2961), .Z(n2946) );
  HDAOI222D2 U3446 ( .A1(n2908), .A2(n3108), .B1(n2866), .B2(n2959), .C1(n3458), .C2(n2906), .Z(n2905) );
  HDAOI22D1 U3447 ( .A1(n2170), .A2(n3071), .B1(n3070), .B2(
        byp_alu_rs1_data_e[20]), .Z(n3073) );
  HDAOI22D1 U3448 ( .A1(n2695), .A2(n3364), .B1(n2682), .B2(n3139), .Z(n2889)
         );
  HDNAN3D1 U3449 ( .A1(n2819), .A2(n3059), .A3(n2961), .Z(n3011) );
  HDNAN3D1 U3450 ( .A1(n2884), .A2(n3107), .A3(n2961), .Z(n3084) );
  HDAND3D1 U3451 ( .A1(n3095), .A2(n2961), .A3(n2868), .Z(n3060) );
  HDNOR2D1 U3452 ( .A1(n2001), .A2(n2456), .Z(n3386) );
  HDAOI22D1 U3453 ( .A1(byp_alu_rs1_data_e[58]), .A2(n2596), .B1(n2597), .B2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_26_), .Z(n2594) );
  HDNAN2D1 U3454 ( .A1(n1767), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_26_), .Z(n2599) );
  HDINVD1 U3455 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_26_), .Z(
        n2600) );
  HDNOR2D1 U3456 ( .A1(n2583), .A2(n3288), .Z(n2584) );
  HDNAN2D1 U3457 ( .A1(n2690), .A2(byp_alu_rs1_data_e[21]), .Z(n2509) );
  HDOAI21M20D1 U3458 ( .A1(byp_alu_rs1_data_e[39]), .A2(n2745), .B(n2677), .Z(
        n3112) );
  HDAND2DL U3459 ( .A1(n3548), .A2(n3549), .Z(n2616) );
  HDNAN2DL U3460 ( .A1(n3556), .A2(ecl_shft_shift4_e[2]), .Z(n3557) );
  HDNAN2D1 U3461 ( .A1(n2698), .A2(byp_alu_rs1_data_e[62]), .Z(n3552) );
  HDOAI211D1 U3462 ( .A1(n3524), .A2(n2710), .B(n3523), .C(n3522), .Z(n3547)
         );
  HDNOR2D1 U3463 ( .A1(n3515), .A2(n2704), .Z(n3516) );
  HDNOR2D2 U3464 ( .A1(n1795), .A2(ecl_shft_lshift_e_l), .Z(n3546) );
  HDNAN2D2 U3465 ( .A1(n2743), .A2(byp_alu_rs1_data_e[10]), .Z(n3513) );
  HDOAI211D1 U3466 ( .A1(n1744), .A2(n3477), .B(n3476), .C(n3475), .Z(n3556)
         );
  HDNOR2D1 U3467 ( .A1(n3472), .A2(n2456), .Z(n3473) );
  HDINVD1 U3468 ( .A(n3364), .Z(n2669) );
  HDAOI22D1 U3469 ( .A1(n3550), .A2(byp_alu_rs1_data_e[20]), .B1(n2653), .B2(
        byp_alu_rs1_data_e[36]), .Z(n3460) );
  HDOAI211D1 U3470 ( .A1(n1743), .A2(n3486), .B(n3485), .C(n3484), .Z(n3570)
         );
  HDNAN2D2 U3471 ( .A1(n2743), .A2(byp_alu_rs1_data_e[9]), .Z(n3505) );
  HDNAN2D2 U3472 ( .A1(n2756), .A2(ecl_alu_log_sel_move_e), .Z(n3278) );
  HDEXOR2D1 U3473 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[36]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_4_) );
  HDAOI211D1 U3474 ( .A1(n1786), .A2(n3008), .B(n2735), .C(n3265), .Z(n2737)
         );
  HDAOI21M20D1 U3475 ( .A1(n3037), .A2(n3561), .B(n2556), .Z(n2558) );
  HDOAI22D1 U3476 ( .A1(n3096), .A2(n3521), .B1(n3565), .B2(n3040), .Z(n3041)
         );
  HDNAN2DL U3477 ( .A1(n1782), .A2(n3112), .Z(n3113) );
  HDAOI21M20D1 U3478 ( .A1(ecl_shft_shift4_e[2]), .A2(ecl_shft_shift4_e[3]), 
        .B(n3575), .Z(n3495) );
  HDAOI211D1 U3479 ( .A1(n2959), .A2(n3474), .B(n2958), .C(n2957), .Z(n3013)
         );
  HDAOI211D1 U3480 ( .A1(n3018), .A2(n3445), .B(n2979), .C(n2978), .Z(n3026)
         );
  HDAOI211D2 U3481 ( .A1(n3298), .A2(ecl_shft_shift4_e[0]), .B(n3087), .C(
        n3086), .Z(n3118) );
  HDOAI22D1 U3482 ( .A1(n3096), .A2(n3505), .B1(n3394), .B2(n3040), .Z(n3006)
         );
  HDOAI22D1 U3483 ( .A1(n3096), .A2(n3498), .B1(n3383), .B2(n3040), .Z(n2997)
         );
  HDAOI211D1 U3484 ( .A1(n2959), .A2(n3464), .B(n2944), .C(n2943), .Z(n2995)
         );
  HDAOI211D2 U3485 ( .A1(ecl_shft_shift4_e[0]), .A2(n3308), .B(n3098), .C(
        n3097), .Z(n3136) );
  HDNOR2D1 U3486 ( .A1(n2675), .A2(n3437), .Z(n3297) );
  HDNAN2D2 U3487 ( .A1(n2743), .A2(byp_alu_rs1_data_e[14]), .Z(n3553) );
  HDAOI22D1 U3488 ( .A1(n1786), .A2(n1756), .B1(n2682), .B2(n3120), .Z(n2884)
         );
  HDAOI21D1 U3489 ( .A1(n2681), .A2(n3258), .B(n2181), .Z(n3002) );
  HDOAI21M20D1 U3490 ( .A1(byp_alu_rs1_data_e[32]), .A2(n2745), .B(n2659), .Z(
        n3008) );
  HDINVDL U3491 ( .A(n2110), .Z(n2533) );
  HDNOR2D2 U3492 ( .A1(n2930), .A2(n2929), .Z(n2982) );
  HDAOI222D2 U3493 ( .A1(n2908), .A2(n2907), .B1(n3445), .B2(n2959), .C1(n3483), .C2(n2906), .Z(n2966) );
  HDAOI222D2 U3494 ( .A1(n2908), .A2(n3143), .B1(n2888), .B2(n2959), .C1(n3474), .C2(n2906), .Z(n2942) );
  HDAOI222D2 U3495 ( .A1(n2908), .A2(n3124), .B1(n2883), .B2(n2959), .C1(n3464), .C2(n2906), .Z(n2924) );
  HDNOR2D2 U3496 ( .A1(n2870), .A2(n2869), .Z(n2904) );
  HDAOI211D2 U3497 ( .A1(n2907), .A2(n1782), .B(n3375), .C(n2722), .Z(n2867)
         );
  HDNOR2D2 U3498 ( .A1(n3116), .A2(n3115), .Z(n3156) );
  HDNOR2D2 U3499 ( .A1(n3122), .A2(n3121), .Z(n3186) );
  HDNOR2D2 U3500 ( .A1(n3162), .A2(n3161), .Z(n3226) );
  HDNOR2D2 U3501 ( .A1(n3064), .A2(n3063), .Z(n3103) );
  HDNOR2D2 U3502 ( .A1(n3004), .A2(n3003), .Z(n3037) );
  HDNOR2D2 U3503 ( .A1(n3181), .A2(n3180), .Z(n3246) );
  HDOAI22D1 U3504 ( .A1(n3469), .A2(n3561), .B1(n3433), .B2(n2702), .Z(n2528)
         );
  HDAOI211D2 U3505 ( .A1(ecl_shft_shift4_e[0]), .A2(n3367), .B(n3366), .C(
        n3365), .Z(n3395) );
  HDOAI21M20D1 U3506 ( .A1(alu_adder_out[40]), .A2(n1785), .B(n2578), .Z(
        alu_byp_rd_data_e[40]) );
  HDOA21M20D2 U3507 ( .A1(n1782), .A2(n3283), .B(n2658), .Z(n3390) );
  HDOA21M20D2 U3508 ( .A1(n1782), .A2(n3295), .B(n2657), .Z(n3399) );
  HDOA21M20D2 U3509 ( .A1(n3318), .A2(n1782), .B(n2658), .Z(n3429) );
  HDOA21M20D2 U3510 ( .A1(n1782), .A2(n3301), .B(n2658), .Z(n3408) );
  HDOA21M20D2 U3511 ( .A1(n1782), .A2(n3327), .B(n2658), .Z(n3434) );
  HDOA21M20D2 U3512 ( .A1(n3336), .A2(n1782), .B(n2657), .Z(n3443) );
  HDAOI21M20D2 U3513 ( .A1(n3521), .A2(n2675), .B(n3163), .Z(n3341) );
  HDOA21M20D2 U3514 ( .A1(n3464), .A2(n2682), .B(n3077), .Z(n3287) );
  HDOA21M20D2 U3515 ( .A1(n3529), .A2(n2680), .B(n3182), .Z(n3349) );
  HDOA21M20D2 U3516 ( .A1(n3458), .A2(n2681), .B(n3059), .Z(n3264) );
  HDOAI21M20D1 U3517 ( .A1(byp_alu_rs1_data_e[43]), .A2(n2745), .B(n2677), .Z(
        n3177) );
  HDNAN2D6 U3518 ( .A1(n1982), .A2(ecl_shft_extendbit_e), .Z(n3260) );
  HDAOI211D2 U3519 ( .A1(ecl_shft_shift4_e[0]), .A2(n3457), .B(n3456), .C(
        n3455), .Z(n3491) );
  HDAOI211D2 U3520 ( .A1(ecl_shft_shift4_e[1]), .A2(n3502), .B(n3495), .C(
        n3463), .Z(n3492) );
  HDAOI211D2 U3521 ( .A1(ecl_shft_shift4_e[1]), .A2(n3510), .B(n3495), .C(
        n3473), .Z(n3501) );
  HDAOI21M20D2 U3522 ( .A1(n1776), .A2(n2669), .B(n3379), .Z(n3472) );
  HDAOI211D2 U3523 ( .A1(ecl_shft_shift4_e[1]), .A2(n3528), .B(n3495), .C(
        n3494), .Z(n3519) );
  HDNAN2D2 U3524 ( .A1(n2743), .A2(byp_alu_rs1_data_e[15]), .Z(n3565) );
  HDAOI211D2 U3525 ( .A1(ecl_shft_shift4_e[1]), .A2(n3520), .B(n3495), .C(
        n3482), .Z(n3509) );
  HDINVDL U3526 ( .A(alu_addsub_rs2_data[17]), .Z(n2572) );
  HDOAI22D1 U3527 ( .A1(n2752), .A2(n2751), .B1(n2766), .B2(n2765), .Z(n2753)
         );
  HDNOR2D2 U3528 ( .A1(n2806), .A2(n2805), .Z(n2848) );
  HDNOR2D2 U3529 ( .A1(n2731), .A2(n2732), .Z(n2785) );
  HDAOI21M20D1 U3530 ( .A1(n2716), .A2(n2456), .B(n2715), .Z(n2721) );
  HDNAN2DL U3531 ( .A1(n1767), .A2(n2131), .Z(n2626) );
  HDAOI21M20D1 U3532 ( .A1(n3157), .A2(n1789), .B(n2630), .Z(n2629) );
  HDAOI211D2 U3533 ( .A1(ecl_shft_shift4_e[0]), .A2(n3373), .B(n3372), .C(
        n3371), .Z(n3397) );
  HDAOI211D2 U3534 ( .A1(ecl_shft_shift4_e[0]), .A2(n3467), .B(n3360), .C(
        n3359), .Z(n3387) );
  HDAOI211D2 U3535 ( .A1(ecl_shft_shift4_e[3]), .A2(n3502), .B(n3392), .C(
        n3391), .Z(n3415) );
  HDOA21M20D2 U3536 ( .A1(n3449), .A2(ecl_shft_shift4_e[0]), .B(n2577), .Z(
        n3368) );
  HDAOI211D2 U3537 ( .A1(ecl_shft_shift4_e[3]), .A2(n3323), .B(n3322), .C(
        n3321), .Z(n3342) );
  HDOR2D1 U3538 ( .A1(n2693), .A2(n3431), .Z(n2504) );
  HDAOI211D2 U3539 ( .A1(ecl_shft_shift4_e[3]), .A2(n3510), .B(n3401), .C(
        n3400), .Z(n3428) );
  HDAOI211D2 U3540 ( .A1(ecl_shft_shift4_e[2]), .A2(n3461), .B(n3424), .C(
        n3423), .Z(n3450) );
  HDAOI211D2 U3541 ( .A1(ecl_shft_shift4_e[3]), .A2(n3449), .B(n2513), .C(
        n2512), .Z(n3470) );
  HDOAI21M20D1 U3542 ( .A1(byp_alu_rs1_data_e[49]), .A2(n2745), .B(n2659), .Z(
        n3295) );
  HDOAI21M20D1 U3543 ( .A1(byp_alu_rs1_data_e[45]), .A2(n2745), .B(n2676), .Z(
        n3216) );
  HDOA21M20D2 U3544 ( .A1(n3445), .A2(n2681), .B(n3039), .Z(n3241) );
  HDOAI21M20D1 U3545 ( .A1(byp_alu_rs1_data_e[38]), .A2(n2745), .B(n2676), .Z(
        n3100) );
  HDNAN2D1 U3546 ( .A1(n1782), .A2(n3237), .Z(n3238) );
  HDOAI21M20D1 U3547 ( .A1(byp_alu_rs1_data_e[46]), .A2(n2745), .B(n2678), .Z(
        n3237) );
  HDOA21M20D2 U3548 ( .A1(n3535), .A2(n2680), .B(n3201), .Z(n3358) );
  HDOAI21M20D1 U3549 ( .A1(byp_alu_rs1_data_e[48]), .A2(n2745), .B(n2676), .Z(
        n3283) );
  HDOAI21M20D1 U3550 ( .A1(byp_alu_rs1_data_e[40]), .A2(n2745), .B(n2676), .Z(
        n3120) );
  HDINVBD4 U3551 ( .A(n1773), .Z(n2681) );
  HDOAI21M20D1 U3552 ( .A1(byp_alu_rs1_data_e[47]), .A2(n2745), .B(n2677), .Z(
        n3258) );
  HDOAI21M20D1 U3553 ( .A1(byp_alu_rs1_data_e[35]), .A2(n2745), .B(n2676), .Z(
        n3061) );
  HDOAI21M20D1 U3554 ( .A1(byp_alu_rs1_data_e[62]), .A2(n2745), .B(n2678), .Z(
        n3407) );
  HDNAN2D8 U3555 ( .A1(n2505), .A2(byp_alu_rs2_data_e[4]), .Z(n3566) );
  HDNAN2D2 U3556 ( .A1(n2712), .A2(ecl_shft_op32_e), .Z(n2744) );
  HDAND2D1 U3557 ( .A1(n2758), .A2(n1769), .Z(n2673) );
  HDAOI211D2 U3558 ( .A1(ecl_shft_shift4_e[0]), .A2(n3084), .B(n3083), .C(
        n3082), .Z(n3105) );
  HDNOR2D2 U3559 ( .A1(n3566), .A2(n3575), .Z(n3001) );
  HDOAI21M20D1 U3560 ( .A1(alu_adder_out[50]), .A2(n1785), .B(n2514), .Z(
        alu_byp_rd_data_e[50]) );
  HDOA211D1 U3561 ( .A1(n2515), .A2(ecl_alu_out_sel_shift_e_l), .B(n2516), .C(
        n2517), .Z(n2514) );
  HDOAI21M20D1 U3562 ( .A1(alu_adder_out[58]), .A2(n1785), .B(n2592), .Z(
        alu_byp_rd_data_e[58]) );
  HDOAI21M20D1 U3563 ( .A1(alu_adder_out[48]), .A2(n1785), .B(n3426), .Z(
        alu_byp_rd_data_e[48]) );
  HDOAI21M20D1 U3564 ( .A1(byp_alu_rs1_data_e[44]), .A2(n2745), .B(n2676), .Z(
        n3196) );
  HDAOI211D1 U3565 ( .A1(n3547), .A2(n3546), .B(n2616), .C(n2617), .Z(n2615)
         );
  HDOAI21M20D1 U3566 ( .A1(n1782), .A2(n3344), .B(n2657), .Z(n3457) );
  HDOAI21M20D1 U3567 ( .A1(byp_alu_rs1_data_e[55]), .A2(n2745), .B(n2676), .Z(
        n3344) );
  HDOAI21M20D1 U3568 ( .A1(n1782), .A2(n3398), .B(n2657), .Z(n3510) );
  HDOAI21M20D1 U3569 ( .A1(byp_alu_rs1_data_e[61]), .A2(n2745), .B(n2659), .Z(
        n3398) );
  HDOAI21M20D1 U3570 ( .A1(n1782), .A2(n3407), .B(n2657), .Z(n3520) );
  HDNOR2D2 U3571 ( .A1(n2158), .A2(ecl_shft_op32_e), .Z(n2505) );
  HDOAI21M20D1 U3572 ( .A1(n1782), .A2(n3389), .B(n2658), .Z(n3502) );
  HDOAI211D1 U3573 ( .A1(n2784), .A2(ecl_alu_out_sel_shift_e_l), .B(n2783), 
        .C(n2782), .Z(alu_byp_rd_data_e[2]) );
  HDOAI21D1 U3574 ( .A1(n2703), .A2(byp_alu_rs1_data_e[2]), .B(n1769), .Z(
        n2781) );
  HDAOI22D1 U3575 ( .A1(byp_alu_rs2_data_e[2]), .A2(n2683), .B1(
        alu_adder_out[2]), .B2(n1785), .Z(n2783) );
  HDOAI211D1 U3576 ( .A1(ecl_alu_out_sel_shift_e_l), .A2(n2816), .B(n2815), 
        .C(n2814), .Z(alu_byp_rd_data_e[4]) );
  HDAOI22D1 U3577 ( .A1(byp_alu_rs2_data_e[4]), .A2(n2683), .B1(
        alu_adder_out[4]), .B2(n1785), .Z(n2814) );
  HDOAI21D1 U3578 ( .A1(n2703), .A2(byp_alu_rs1_data_e[4]), .B(n1769), .Z(
        n2813) );
  HDNOR4D1 U3579 ( .A1(n2811), .A2(n2810), .A3(n2809), .A4(n2808), .Z(n2816)
         );
  HDOAI22D1 U3580 ( .A1(n2807), .A2(n2686), .B1(n2836), .B2(n3560), .Z(n2808)
         );
  HDOAI22D1 U3581 ( .A1(n2849), .A2(n1789), .B1(n2848), .B2(n3561), .Z(n2810)
         );
  HDOAI22D1 U3582 ( .A1(n2837), .A2(n3563), .B1(n2802), .B2(n2702), .Z(n2811)
         );
  HDOAI211D1 U3583 ( .A1(ecl_alu_out_sel_shift_e_l), .A2(n2801), .B(n2800), 
        .C(n2799), .Z(alu_byp_rd_data_e[3]) );
  HDOAI21D1 U3584 ( .A1(n2703), .A2(byp_alu_rs1_data_e[3]), .B(n1769), .Z(
        n2798) );
  HDNOR4D1 U3585 ( .A1(n2796), .A2(n2795), .A3(n2794), .A4(n2793), .Z(n2801)
         );
  HDOAI22D1 U3586 ( .A1(n2792), .A2(n2686), .B1(n2836), .B2(n3561), .Z(n2793)
         );
  HDOAI22D1 U3587 ( .A1(n1789), .A2(n2837), .B1(n2802), .B2(n3576), .Z(n2795)
         );
  HDOAI211D1 U3588 ( .A1(n2561), .A2(n2562), .B(n2563), .C(n2564), .Z(
        alu_byp_rd_data_e[17]) );
  HDNOR4D1 U3589 ( .A1(n2567), .A2(n2566), .A3(n2568), .A4(n2565), .Z(n2561)
         );
  HDAOI22D1 U3590 ( .A1(byp_alu_rs2_data_e[17]), .A2(n2683), .B1(n2571), .B2(
        byp_alu_rs1_data_e[17]), .Z(n2570) );
  HDOAI21D1 U3591 ( .A1(n2703), .A2(byp_alu_rs1_data_e[17]), .B(n1769), .Z(
        n2569) );
  HDOAI22D1 U3592 ( .A1(n3013), .A2(n2686), .B1(n3038), .B2(n3563), .Z(n2568)
         );
  HDOAI22D1 U3593 ( .A1(n3012), .A2(n2702), .B1(n3057), .B2(n3561), .Z(n2567)
         );
  HDAO21M20D1 U3594 ( .A1(n3037), .A2(n3560), .B(n2573), .Z(n2566) );
  HDAOI22D1 U3595 ( .A1(byp_alu_rs2_data_e[6]), .A2(n2683), .B1(
        alu_adder_out[6]), .B2(n1785), .Z(n2845) );
  HDNAN2D1 U3596 ( .A1(n2842), .A2(n1769), .Z(n2843) );
  HDOAI21D1 U3597 ( .A1(n2703), .A2(byp_alu_rs1_data_e[6]), .B(n1769), .Z(
        n2844) );
  HDNOR4D1 U3598 ( .A1(n2840), .A2(n2841), .A3(n2839), .A4(n2838), .Z(n2847)
         );
  HDOAI22D1 U3599 ( .A1(n2837), .A2(n2686), .B1(n2836), .B2(n2702), .Z(n2838)
         );
  HDOAI22D1 U3600 ( .A1(n2882), .A2(n1789), .B1(n2881), .B2(n3561), .Z(n2839)
         );
  HDOAI22D1 U3601 ( .A1(n2865), .A2(n3563), .B1(n2864), .B2(n3560), .Z(n2840)
         );
  HDOAI22D1 U3602 ( .A1(n2849), .A2(n1783), .B1(n2848), .B2(n3576), .Z(n2841)
         );
  HDAOI22D1 U3603 ( .A1(n1742), .A2(n2683), .B1(alu_adder_out[5]), .B2(n1785), 
        .Z(n2829) );
  HDNAN2D1 U3604 ( .A1(n2826), .A2(n1769), .Z(n2827) );
  HDOAI21D1 U3605 ( .A1(n2703), .A2(byp_alu_rs1_data_e[5]), .B(n1769), .Z(
        n2828) );
  HDOAI22D1 U3606 ( .A1(n2822), .A2(n2686), .B1(n2836), .B2(n3576), .Z(n2823)
         );
  HDAOI22D1 U3607 ( .A1(n2789), .A2(ecl_shft_shift4_e[0]), .B1(n2850), .B2(
        ecl_shft_shift4_e[1]), .Z(n2790) );
  HDNAN2D1 U3608 ( .A1(n2981), .A2(ecl_shft_shift4_e[3]), .Z(n2791) );
  HDOAI22D1 U3609 ( .A1(n2865), .A2(n1789), .B1(n2455), .B2(n3561), .Z(n2824)
         );
  HDOAI22D1 U3610 ( .A1(n2849), .A2(n3563), .B1(n2848), .B2(n3560), .Z(n2825)
         );
  HDAOI22D1 U3611 ( .A1(n2962), .A2(ecl_shft_shift4_e[3]), .B1(
        ecl_shft_shift4_e[1]), .B2(n2832), .Z(n2777) );
  HDAOI22D1 U3612 ( .A1(byp_alu_rs2_data_e[15]), .A2(n2683), .B1(
        alu_adder_out[15]), .B2(n1785), .Z(n2991) );
  HDAOI22D1 U3613 ( .A1(n2145), .A2(n2990), .B1(n2989), .B2(
        byp_alu_rs1_data_e[15]), .Z(n2992) );
  HDNAN2D1 U3614 ( .A1(n2988), .A2(n1769), .Z(n2989) );
  HDOAI21D1 U3615 ( .A1(n2703), .A2(byp_alu_rs1_data_e[15]), .B(n1769), .Z(
        n2990) );
  HDNOR4D1 U3616 ( .A1(n2987), .A2(n2986), .A3(n2985), .A4(n2984), .Z(n2993)
         );
  HDOAI22D1 U3617 ( .A1(n2983), .A2(n2686), .B1(n2982), .B2(n2702), .Z(n2984)
         );
  HDOAI22D1 U3618 ( .A1(n3026), .A2(n1789), .B1(n3025), .B2(n3561), .Z(n2985)
         );
  HDOAI22D1 U3619 ( .A1(n3013), .A2(n3563), .B1(n3012), .B2(n3560), .Z(n2986)
         );
  HDOAI22D1 U3620 ( .A1(n2995), .A2(n1783), .B1(n2994), .B2(n3576), .Z(n2987)
         );
  HDNAN4D1 U3621 ( .A1(n2634), .A2(n2632), .A3(n2633), .A4(n2631), .Z(
        alu_byp_rd_data_e[21]) );
  HDNAN2D1 U3622 ( .A1(alu_adder_out[21]), .A2(n1785), .Z(n2631) );
  HDOR2D1 U3623 ( .A1(n3105), .A2(n2642), .Z(n2633) );
  HDOR2D1 U3624 ( .A1(n3561), .A2(ecl_alu_out_sel_shift_e_l), .Z(n2642) );
  HDNOR2D1 U3625 ( .A1(n2638), .A2(n2639), .Z(n2632) );
  HDNOR3D1 U3626 ( .A1(n3093), .A2(ecl_alu_out_sel_shift_e_l), .A3(n3576), .Z(
        n2638) );
  HDOAI31D1 U3627 ( .A1(n2635), .A2(n2636), .A3(n2637), .B(n1924), .Z(n2634)
         );
  HDOAI222D1 U3628 ( .A1(n3094), .A2(n1783), .B1(n3106), .B2(n1789), .C1(n3104), .C2(n3563), .Z(n2637) );
  HDNOR2D1 U3629 ( .A1(n3103), .A2(n3560), .Z(n2636) );
  HDOAI22D1 U3630 ( .A1(n3075), .A2(n2702), .B1(n3076), .B2(n3533), .Z(n2635)
         );
  HDAOI21D1 U3631 ( .A1(alu_adder_out[9]), .A2(n1785), .B(n2539), .Z(n2538) );
  HDAOI22D1 U3632 ( .A1(byp_alu_rs2_data_e[8]), .A2(n2683), .B1(
        alu_adder_out[8]), .B2(n1785), .Z(n2878) );
  HDNAN2D1 U3633 ( .A1(n2875), .A2(n1769), .Z(n2876) );
  HDOAI21D1 U3634 ( .A1(n2703), .A2(byp_alu_rs1_data_e[8]), .B(n1769), .Z(
        n2877) );
  HDNOR4D1 U3635 ( .A1(n2874), .A2(n2873), .A3(n2872), .A4(n2871), .Z(n2880)
         );
  HDOAI22D1 U3636 ( .A1(n2894), .A2(n3563), .B1(n2893), .B2(n3560), .Z(n2871)
         );
  HDOAI22D1 U3637 ( .A1(n2882), .A2(n1783), .B1(n2881), .B2(n3576), .Z(n2872)
         );
  HDOAI22D1 U3638 ( .A1(n2905), .A2(n1789), .B1(n2904), .B2(n3561), .Z(n2873)
         );
  HDOAI22D1 U3639 ( .A1(n2865), .A2(n2686), .B1(n2455), .B2(n2702), .Z(n2874)
         );
  HDAOI211D1 U3640 ( .A1(ecl_shft_shift4_e[1]), .A2(n2760), .B(n2739), .C(
        n2738), .Z(n2752) );
  HDOAI211D1 U3641 ( .A1(n2737), .A2(n2456), .B(n2792), .C(n2736), .Z(n2738)
         );
  HDNOR2D1 U3642 ( .A1(n2887), .A2(n2710), .Z(n2739) );
  HDAO21D1 U3643 ( .A1(ecl_shft_shift1_e[2]), .A2(n2764), .B(n2754), .Z(n2666)
         );
  HDAOI22D1 U3644 ( .A1(byp_alu_rs2_data_e[10]), .A2(n2683), .B1(
        alu_adder_out[10]), .B2(n1785), .Z(n2901) );
  HDOAI21D1 U3645 ( .A1(n2703), .A2(byp_alu_rs1_data_e[10]), .B(n1769), .Z(
        n2900) );
  HDNOR4D1 U3646 ( .A1(n2897), .A2(n2898), .A3(n2896), .A4(n2895), .Z(n2903)
         );
  HDOAI22D1 U3647 ( .A1(n2894), .A2(n2686), .B1(n2893), .B2(n2702), .Z(n2895)
         );
  HDOAI22D1 U3648 ( .A1(n2942), .A2(n1789), .B1(n2941), .B2(n3561), .Z(n2896)
         );
  HDOAI22D1 U3649 ( .A1(n2924), .A2(n3563), .B1(n2923), .B2(n3560), .Z(n2897)
         );
  HDOAI22D1 U3650 ( .A1(n2905), .A2(n1783), .B1(n2904), .B2(n3576), .Z(n2898)
         );
  HDAOI22D1 U3651 ( .A1(byp_alu_rs2_data_e[7]), .A2(n2683), .B1(
        alu_adder_out[7]), .B2(n1785), .Z(n2861) );
  HDNAN2D1 U3652 ( .A1(n2858), .A2(n1769), .Z(n2859) );
  HDOAI21D1 U3653 ( .A1(n2703), .A2(byp_alu_rs1_data_e[7]), .B(n1769), .Z(
        n2860) );
  HDNOR4D1 U3654 ( .A1(n2856), .A2(n2857), .A3(n2855), .A4(n2854), .Z(n2863)
         );
  HDOAI22D1 U3655 ( .A1(n2894), .A2(n1789), .B1(n2893), .B2(n3561), .Z(n2854)
         );
  HDAOI22D1 U3656 ( .A1(n3043), .A2(ecl_shft_shift4_e[3]), .B1(n2981), .B2(
        ecl_shft_shift4_e[2]), .Z(n2852) );
  HDNAN2D1 U3657 ( .A1(n2850), .A2(ecl_shft_shift4_e[0]), .Z(n2853) );
  HDAOI22D1 U3658 ( .A1(n2908), .A2(n3483), .B1(n3445), .B2(n2906), .Z(n2894)
         );
  HDOAI22D1 U3659 ( .A1(n2882), .A2(n3563), .B1(n2881), .B2(n3560), .Z(n2855)
         );
  HDAOI22D1 U3660 ( .A1(n2962), .A2(ecl_shft_shift4_e[2]), .B1(
        ecl_shft_shift4_e[3]), .B2(n3022), .Z(n2834) );
  HDAOI22D1 U3661 ( .A1(n2908), .A2(n3474), .B1(n2888), .B2(n2906), .Z(n2882)
         );
  HDOAI22D1 U3662 ( .A1(n2865), .A2(n1783), .B1(n2864), .B2(n3576), .Z(n2856)
         );
  HDNAN2D1 U3663 ( .A1(n2818), .A2(ecl_shft_shift4_e[0]), .Z(n2821) );
  HDAOI22D1 U3664 ( .A1(n2908), .A2(n3464), .B1(n2883), .B2(n2906), .Z(n2865)
         );
  HDOAI22D1 U3665 ( .A1(n2849), .A2(n2686), .B1(n2848), .B2(n2702), .Z(n2857)
         );
  HDOAI22D1 U3666 ( .A1(n2928), .A2(n2709), .B1(n2804), .B2(n2456), .Z(n2805)
         );
  HDOAI22D1 U3667 ( .A1(n2999), .A2(n2710), .B1(n2867), .B2(n2704), .Z(n2806)
         );
  HDAOI22D1 U3668 ( .A1(n2908), .A2(n3458), .B1(n2866), .B2(n2906), .Z(n2849)
         );
  HDOAI211D1 U3669 ( .A1(n3174), .A2(ecl_alu_out_sel_shift_e_l), .B(n3173), 
        .C(n3172), .Z(alu_byp_rd_data_e[27]) );
  HDNAN2D1 U3670 ( .A1(n3169), .A2(n1769), .Z(n3170) );
  HDOAI21D1 U3671 ( .A1(n2703), .A2(byp_alu_rs1_data_e[27]), .B(n1769), .Z(
        n3171) );
  HDOAI22D1 U3672 ( .A1(n3186), .A2(n3576), .B1(n3185), .B2(n1783), .Z(n3167)
         );
  HDOAI22D1 U3673 ( .A1(n3226), .A2(n3561), .B1(n3225), .B2(n1789), .Z(n3168)
         );
  HDOAI211D1 U3674 ( .A1(n3134), .A2(ecl_alu_out_sel_shift_e_l), .B(n3133), 
        .C(n3132), .Z(alu_byp_rd_data_e[25]) );
  HDAOI22D1 U3675 ( .A1(byp_alu_rs2_data_e[25]), .A2(n2683), .B1(
        alu_adder_out[25]), .B2(n1785), .Z(n3132) );
  HDNAN2D1 U3676 ( .A1(n3129), .A2(n1769), .Z(n3130) );
  HDOAI21D1 U3677 ( .A1(n2703), .A2(byp_alu_rs1_data_e[25]), .B(n1769), .Z(
        n3131) );
  HDNOR4D1 U3678 ( .A1(n3128), .A2(n3127), .A3(n3126), .A4(n3125), .Z(n3134)
         );
  HDOAI22D1 U3679 ( .A1(n3186), .A2(n3561), .B1(n3185), .B2(n1789), .Z(n3125)
         );
  HDOAI22D1 U3680 ( .A1(n3136), .A2(n1783), .B1(n3135), .B2(n3576), .Z(n3126)
         );
  HDOAI22D1 U3681 ( .A1(n3157), .A2(n3563), .B1(n2115), .B2(n3560), .Z(n3127)
         );
  HDOAI22D1 U3682 ( .A1(n3118), .A2(n3533), .B1(n3117), .B2(n2702), .Z(n3128)
         );
  HDOAI22D1 U3683 ( .A1(n3105), .A2(n3576), .B1(n3117), .B2(n3560), .Z(n2530)
         );
  HDOA21M20D1 U3684 ( .A1(alu_adder_out[23]), .A2(n1785), .B(n2537), .Z(n2529)
         );
  HDOAI21D1 U3685 ( .A1(n2703), .A2(byp_alu_rs1_data_e[23]), .B(n1769), .Z(
        n2531) );
  HDOAI222D1 U3686 ( .A1(n3104), .A2(n3533), .B1(n3106), .B2(n1783), .C1(n3103), .C2(n2702), .Z(n2536) );
  HDOAI22D1 U3687 ( .A1(n3118), .A2(n3563), .B1(n3135), .B2(n3561), .Z(n2534)
         );
  HDOAI21D1 U3688 ( .A1(n2551), .A2(ecl_alu_out_sel_shift_e_l), .B(n2552), .Z(
        alu_byp_rd_data_e[16]) );
  HDAOI21D1 U3689 ( .A1(alu_adder_out[16]), .A2(n1785), .B(n2553), .Z(n2552)
         );
  HDAND4D1 U3690 ( .A1(n2560), .A2(n2557), .A3(n2558), .A4(n2559), .Z(n2551)
         );
  HDOR2D1 U3691 ( .A1(n2994), .A2(n2702), .Z(n2559) );
  HDOA222D1 U3692 ( .A1(n3012), .A2(n3576), .B1(n3038), .B2(n1789), .C1(n2995), 
        .C2(n2686), .Z(n2557) );
  HDNAN2M1D1 U3693 ( .A1(n3025), .A2(n2692), .Z(n2560) );
  HDAOI22D1 U3694 ( .A1(byp_alu_rs2_data_e[13]), .A2(n2683), .B1(
        alu_adder_out[13]), .B2(n1785), .Z(n2954) );
  HDNAN2D1 U3695 ( .A1(n2951), .A2(n1769), .Z(n2952) );
  HDOAI21D1 U3696 ( .A1(n2703), .A2(byp_alu_rs1_data_e[13]), .B(n1769), .Z(
        n2953) );
  HDNOR4D1 U3697 ( .A1(n2949), .A2(n2950), .A3(n2948), .A4(n2947), .Z(n2956)
         );
  HDOAI22D1 U3698 ( .A1(n2983), .A2(n3563), .B1(n2982), .B2(n3560), .Z(n2947)
         );
  HDOAI22D1 U3699 ( .A1(n2966), .A2(n1783), .B1(n2965), .B2(n3576), .Z(n2948)
         );
  HDOAI22D1 U3700 ( .A1(n2995), .A2(n1789), .B1(n2994), .B2(n3561), .Z(n2949)
         );
  HDOAI22D1 U3701 ( .A1(n2942), .A2(n2686), .B1(n2941), .B2(n2702), .Z(n2950)
         );
  HDOAI211D1 U3702 ( .A1(n2773), .A2(ecl_alu_out_sel_shift_e_l), .B(n2772), 
        .C(n2771), .Z(alu_byp_rd_data_e[1]) );
  HDNAN2D1 U3703 ( .A1(n2768), .A2(n1769), .Z(n2769) );
  HDOAI21D1 U3704 ( .A1(n2703), .A2(byp_alu_rs1_data_e[1]), .B(n1769), .Z(
        n2770) );
  HDAOI22D1 U3705 ( .A1(byp_alu_rs2_data_e[1]), .A2(n2683), .B1(
        alu_adder_out[1]), .B2(n1785), .Z(n2772) );
  HDOAI211D1 U3706 ( .A1(n2867), .A2(n2705), .B(n2726), .C(n2837), .Z(n2732)
         );
  HDNAN2D1 U3707 ( .A1(n2724), .A2(ecl_shft_shift4_e[0]), .Z(n2726) );
  HDOAI211D1 U3708 ( .A1(n2748), .A2(n2456), .B(n2807), .C(n2747), .Z(n2749)
         );
  HDNOR2D1 U3709 ( .A1(n2892), .A2(n2710), .Z(n2750) );
  HDOAI211D1 U3710 ( .A1(n3320), .A2(n2685), .B(n2143), .C(n2740), .Z(n2775)
         );
  HDINVD1 U3711 ( .A(n2764), .Z(n2774) );
  HDOAI211D1 U3712 ( .A1(n2912), .A2(n2710), .B(n2721), .C(n2720), .Z(n2764)
         );
  HDAOI22D1 U3713 ( .A1(n2789), .A2(ecl_shft_shift4_e[1]), .B1(n2850), .B2(
        ecl_shft_shift4_e[2]), .Z(n2720) );
  HDOAI211D1 U3714 ( .A1(n3513), .A2(n2685), .B(n3362), .C(n2719), .Z(n2850)
         );
  HDOAI211D1 U3715 ( .A1(n3331), .A2(n2685), .B(n2507), .C(n2718), .Z(n2789)
         );
  HDAOI211D1 U3716 ( .A1(n3536), .A2(n3301), .B(n3297), .C(n2714), .Z(n2716)
         );
  HDAOI22D1 U3717 ( .A1(n2818), .A2(ecl_shft_shift4_e[1]), .B1(n2946), .B2(
        ecl_shft_shift4_e[3]), .Z(n2762) );
  HDOAI211D1 U3718 ( .A1(n3316), .A2(n2685), .B(n2733), .C(n3315), .Z(n2760)
         );
  HDAOI22D1 U3719 ( .A1(byp_alu_rs2_data_e[12]), .A2(n2683), .B1(
        alu_adder_out[12]), .B2(n1785), .Z(n2938) );
  HDNAN2D1 U3720 ( .A1(n2935), .A2(n1769), .Z(n2936) );
  HDOAI21D1 U3721 ( .A1(n2703), .A2(byp_alu_rs1_data_e[12]), .B(n1769), .Z(
        n2937) );
  HDNOR4D1 U3722 ( .A1(n2934), .A2(n2933), .A3(n2932), .A4(n2931), .Z(n2940)
         );
  HDOAI22D1 U3723 ( .A1(n2983), .A2(n1789), .B1(n2982), .B2(n3561), .Z(n2931)
         );
  HDOAI22D1 U3724 ( .A1(n2966), .A2(n3563), .B1(n2965), .B2(n3560), .Z(n2932)
         );
  HDOAI22D1 U3725 ( .A1(n2942), .A2(n1783), .B1(n2941), .B2(n3576), .Z(n2933)
         );
  HDOAI22D1 U3726 ( .A1(n2924), .A2(n2686), .B1(n2923), .B2(n2702), .Z(n2934)
         );
  HDOAI211D1 U3727 ( .A1(ecl_alu_out_sel_shift_e_l), .A2(n2976), .B(n2975), 
        .C(n2974), .Z(alu_byp_rd_data_e[14]) );
  HDAOI22D1 U3728 ( .A1(byp_alu_rs2_data_e[14]), .A2(n2683), .B1(
        alu_adder_out[14]), .B2(n1785), .Z(n2974) );
  HDNAN2D1 U3729 ( .A1(n2971), .A2(n1769), .Z(n2972) );
  HDOAI21D1 U3730 ( .A1(n2703), .A2(byp_alu_rs1_data_e[14]), .B(n1769), .Z(
        n2973) );
  HDNOR4D1 U3731 ( .A1(n2970), .A2(n2969), .A3(n2968), .A4(n2967), .Z(n2976)
         );
  HDOAI22D1 U3732 ( .A1(n2983), .A2(n1783), .B1(n2982), .B2(n3576), .Z(n2967)
         );
  HDOAI22D1 U3733 ( .A1(n2928), .A2(n2456), .B1(n2999), .B2(n2704), .Z(n2929)
         );
  HDOAI22D1 U3734 ( .A1(n3060), .A2(n2709), .B1(n3111), .B2(n2710), .Z(n2930)
         );
  HDNOR2D1 U3735 ( .A1(n3165), .A2(n3422), .Z(n2926) );
  HDOAI22D1 U3736 ( .A1(n2966), .A2(n2686), .B1(n2965), .B2(n2702), .Z(n2968)
         );
  HDOAI22D1 U3737 ( .A1(n3013), .A2(n1789), .B1(n3012), .B2(n3561), .Z(n2969)
         );
  HDAOI22D1 U3738 ( .A1(n2962), .A2(ecl_shft_shift4_e[0]), .B1(
        ecl_shft_shift4_e[1]), .B2(n3022), .Z(n2963) );
  HDNAN2D1 U3739 ( .A1(n3092), .A2(ecl_shft_shift4_e[2]), .Z(n2964) );
  HDNOR2D1 U3740 ( .A1(n3165), .A2(n3436), .Z(n2958) );
  HDOAI22D1 U3741 ( .A1(n2995), .A2(n3563), .B1(n2994), .B2(n3560), .Z(n2970)
         );
  HDNOR2D1 U3742 ( .A1(n3165), .A2(n3431), .Z(n2944) );
  HDAOI22D1 U3743 ( .A1(byp_alu_rs2_data_e[11]), .A2(n2683), .B1(
        alu_adder_out[11]), .B2(n1785), .Z(n2920) );
  HDNAN2D1 U3744 ( .A1(n2917), .A2(n1769), .Z(n2918) );
  HDOAI21D1 U3745 ( .A1(n2703), .A2(byp_alu_rs1_data_e[11]), .B(n1769), .Z(
        n2919) );
  HDNOR4D1 U3746 ( .A1(n2915), .A2(n2916), .A3(n2914), .A4(n2913), .Z(n2922)
         );
  HDOAI22D1 U3747 ( .A1(n2966), .A2(n1789), .B1(n2965), .B2(n3561), .Z(n2913)
         );
  HDAOI22D1 U3748 ( .A1(n3099), .A2(ecl_shft_shift4_e[3]), .B1(n3043), .B2(
        ecl_shft_shift4_e[2]), .Z(n2910) );
  HDNAN2D1 U3749 ( .A1(n2981), .A2(ecl_shft_shift4_e[1]), .Z(n2911) );
  HDOAI22D1 U3750 ( .A1(n2942), .A2(n3563), .B1(n2941), .B2(n3560), .Z(n2914)
         );
  HDAOI22D1 U3751 ( .A1(n3092), .A2(ecl_shft_shift4_e[3]), .B1(
        ecl_shft_shift4_e[2]), .B2(n3022), .Z(n2890) );
  HDNAN2D1 U3752 ( .A1(n2962), .A2(ecl_shft_shift4_e[1]), .Z(n2891) );
  HDNAN2D1 U3753 ( .A1(n2946), .A2(ecl_shft_shift4_e[1]), .Z(n2886) );
  HDAOI22D1 U3754 ( .A1(n2695), .A2(n3283), .B1(n2680), .B2(n3008), .Z(n2761)
         );
  HDAOI22D1 U3755 ( .A1(n1786), .A2(n3196), .B1(n3536), .B2(n3389), .Z(n2734)
         );
  HDOAI22D1 U3756 ( .A1(n2905), .A2(n2686), .B1(n2904), .B2(n2702), .Z(n2916)
         );
  HDOAI22D1 U3757 ( .A1(n3060), .A2(n2710), .B1(n2999), .B2(n2707), .Z(n2869)
         );
  HDOAI22D1 U3758 ( .A1(n2928), .A2(n2704), .B1(n2867), .B2(n2456), .Z(n2870)
         );
  HDOAI22M10D1 U3759 ( .A1(n3177), .A2(n2654), .B1(n3175), .B2(n3566), .Z(
        n2722) );
  HDAOI22D1 U3760 ( .A1(n2727), .A2(n1782), .B1(n3418), .B2(n3536), .Z(n2728)
         );
  HDINVD1 U3761 ( .A(n3565), .Z(n2727) );
  HDOAI211D1 U3762 ( .A1(ecl_alu_out_sel_shift_e_l), .A2(n3036), .B(n3035), 
        .C(n3034), .Z(alu_byp_rd_data_e[18]) );
  HDAOI22D1 U3763 ( .A1(byp_alu_rs2_data_e[18]), .A2(n2683), .B1(
        alu_adder_out[18]), .B2(n1785), .Z(n3034) );
  HDNAN2D1 U3764 ( .A1(n3031), .A2(n1769), .Z(n3032) );
  HDOAI21D1 U3765 ( .A1(n2703), .A2(byp_alu_rs1_data_e[18]), .B(n1769), .Z(
        n3033) );
  HDNOR4D1 U3766 ( .A1(n3030), .A2(n3029), .A3(n3028), .A4(n3027), .Z(n3036)
         );
  HDOAI22D1 U3767 ( .A1(n2453), .A2(n2686), .B1(n3025), .B2(n2702), .Z(n3027)
         );
  HDINVD1 U3768 ( .A(n3044), .Z(n2788) );
  HDNOR2D1 U3769 ( .A1(n3096), .A2(n3340), .Z(n2979) );
  HDOAI22D1 U3770 ( .A1(n3038), .A2(n1783), .B1(n3037), .B2(n3576), .Z(n3028)
         );
  HDOAI22D1 U3771 ( .A1(n3076), .A2(n1789), .B1(n3075), .B2(n3561), .Z(n3029)
         );
  HDOAI22D1 U3772 ( .A1(n3058), .A2(n3563), .B1(n3057), .B2(n3560), .Z(n3030)
         );
  HDOAI211D1 U3773 ( .A1(n2620), .A2(ecl_alu_out_sel_shift_e_l), .B(n2621), 
        .C(n2622), .Z(alu_byp_rd_data_e[24]) );
  HDOAI22D1 U3774 ( .A1(n3576), .A2(n3117), .B1(n3105), .B2(n2702), .Z(n2623)
         );
  HDAOI21D1 U3775 ( .A1(alu_adder_out[24]), .A2(n1785), .B(n2624), .Z(n2621)
         );
  HDNOR2D1 U3776 ( .A1(n2627), .A2(n2628), .Z(n2620) );
  HDOAI21D1 U3777 ( .A1(n3135), .A2(n3560), .B(n2629), .Z(n2628) );
  HDOAI22D1 U3778 ( .A1(n3106), .A2(n3533), .B1(n3156), .B2(n3561), .Z(n2630)
         );
  HDOAI22D1 U3779 ( .A1(n3118), .A2(n1783), .B1(n3136), .B2(n3563), .Z(n2627)
         );
  HDOAI211D1 U3780 ( .A1(n3215), .A2(ecl_alu_out_sel_shift_e_l), .B(n3214), 
        .C(n3213), .Z(alu_byp_rd_data_e[29]) );
  HDAOI22D1 U3781 ( .A1(byp_alu_rs2_data_e[29]), .A2(n2683), .B1(
        alu_adder_out[29]), .B2(n1785), .Z(n3213) );
  HDNAN2D1 U3782 ( .A1(n3210), .A2(n1769), .Z(n3211) );
  HDOAI21D1 U3783 ( .A1(n2703), .A2(byp_alu_rs1_data_e[29]), .B(n1769), .Z(
        n3212) );
  HDNOR4D1 U3784 ( .A1(n3206), .A2(n3208), .A3(n3207), .A4(n3209), .Z(n3215)
         );
  HDOAI22D1 U3785 ( .A1(n3226), .A2(n3576), .B1(n3225), .B2(n1783), .Z(n3207)
         );
  HDOAI22D1 U3786 ( .A1(n3246), .A2(n3560), .B1(n3245), .B2(n3563), .Z(n3209)
         );
  HDOAI211D1 U3787 ( .A1(ecl_alu_out_sel_shift_e_l), .A2(n3236), .B(n3235), 
        .C(n3234), .Z(alu_byp_rd_data_e[30]) );
  HDAOI22D1 U3788 ( .A1(byp_alu_rs2_data_e[30]), .A2(n2683), .B1(
        alu_adder_out[30]), .B2(n1785), .Z(n3234) );
  HDNAN2D1 U3789 ( .A1(n3231), .A2(n1769), .Z(n3232) );
  HDOAI21D1 U3790 ( .A1(n2703), .A2(byp_alu_rs1_data_e[30]), .B(n1769), .Z(
        n3233) );
  HDNOR4D1 U3791 ( .A1(n3230), .A2(n3229), .A3(n3228), .A4(n3227), .Z(n3236)
         );
  HDOAI22D1 U3792 ( .A1(n3226), .A2(n2702), .B1(n3225), .B2(n3533), .Z(n3227)
         );
  HDOAI22D1 U3793 ( .A1(n3292), .A2(n3561), .B1(n3291), .B2(n1789), .Z(n3228)
         );
  HDOAI22D1 U3794 ( .A1(n3246), .A2(n3576), .B1(n3245), .B2(n1783), .Z(n3230)
         );
  HDOAI211D1 U3795 ( .A1(ecl_alu_out_sel_shift_e_l), .A2(n3155), .B(n3154), 
        .C(n3153), .Z(alu_byp_rd_data_e[26]) );
  HDAOI22D1 U3796 ( .A1(byp_alu_rs2_data_e[26]), .A2(n2683), .B1(
        alu_adder_out[26]), .B2(n1785), .Z(n3153) );
  HDNAN2D1 U3797 ( .A1(n3150), .A2(n1769), .Z(n3151) );
  HDOAI21D1 U3798 ( .A1(n2703), .A2(byp_alu_rs1_data_e[26]), .B(n1769), .Z(
        n3152) );
  HDNOR4D1 U3799 ( .A1(n3149), .A2(n3148), .A3(n3147), .A4(n3146), .Z(n3155)
         );
  HDOAI22D1 U3800 ( .A1(n3186), .A2(n3560), .B1(n3185), .B2(n3563), .Z(n3147)
         );
  HDOAI22D1 U3801 ( .A1(n3136), .A2(n3533), .B1(n3135), .B2(n2702), .Z(n3148)
         );
  HDNAN2D1 U3802 ( .A1(n3099), .A2(ecl_shft_shift4_e[0]), .Z(n3102) );
  HDNOR2D1 U3803 ( .A1(n3241), .A2(n2704), .Z(n3097) );
  HDOAI22D1 U3804 ( .A1(n3165), .A2(n3521), .B1(n3565), .B2(n3096), .Z(n3098)
         );
  HDOAI22D1 U3805 ( .A1(n3157), .A2(n1783), .B1(n2115), .B2(n3576), .Z(n3149)
         );
  HDOAI22D1 U3806 ( .A1(n3383), .A2(n3165), .B1(n3184), .B2(n2707), .Z(n3109)
         );
  HDOAI22D1 U3807 ( .A1(n3264), .A2(n2704), .B1(n3183), .B2(n2456), .Z(n3110)
         );
  HDOAI211D1 U3808 ( .A1(ecl_alu_out_sel_shift_e_l), .A2(n3195), .B(n3194), 
        .C(n3193), .Z(alu_byp_rd_data_e[28]) );
  HDAOI22D1 U3809 ( .A1(byp_alu_rs2_data_e[28]), .A2(n2683), .B1(
        alu_adder_out[28]), .B2(n1785), .Z(n3193) );
  HDNAN2D1 U3810 ( .A1(n3190), .A2(n1769), .Z(n3191) );
  HDOAI21D1 U3811 ( .A1(n2703), .A2(byp_alu_rs1_data_e[28]), .B(n1769), .Z(
        n3192) );
  HDNOR2D1 U3812 ( .A1(n3332), .A2(n2456), .Z(n3144) );
  HDOAI22D1 U3813 ( .A1(n3553), .A2(n3165), .B1(n3224), .B2(n2705), .Z(n3145)
         );
  HDOAI22D1 U3814 ( .A1(n3296), .A2(n2708), .B1(n3328), .B2(n2710), .Z(n3140)
         );
  HDOAI22D1 U3815 ( .A1(n3220), .A2(n2704), .B1(n3137), .B2(n2456), .Z(n3141)
         );
  HDOAI22D1 U3816 ( .A1(n3186), .A2(n2702), .B1(n3185), .B2(n3533), .Z(n3188)
         );
  HDOAI22D1 U3817 ( .A1(n3284), .A2(n2709), .B1(n3319), .B2(n2710), .Z(n3121)
         );
  HDOAI22D1 U3818 ( .A1(n3200), .A2(n2704), .B1(n3119), .B2(n2456), .Z(n3122)
         );
  HDOAI22D1 U3819 ( .A1(n3335), .A2(n2710), .B1(n3302), .B2(n2708), .Z(n3161)
         );
  HDOAI22D1 U3820 ( .A1(n3240), .A2(n2704), .B1(n3158), .B2(n2456), .Z(n3162)
         );
  HDOAI211D1 U3821 ( .A1(ecl_alu_out_sel_shift_e_l), .A2(n3074), .B(n3073), 
        .C(n3072), .Z(alu_byp_rd_data_e[20]) );
  HDAOI22D1 U3822 ( .A1(byp_alu_rs2_data_e[20]), .A2(n2683), .B1(
        alu_adder_out[20]), .B2(n1785), .Z(n3072) );
  HDNAN2D1 U3823 ( .A1(n3069), .A2(n1769), .Z(n3070) );
  HDOAI21D1 U3824 ( .A1(n2703), .A2(byp_alu_rs1_data_e[20]), .B(n1769), .Z(
        n3071) );
  HDNOR4D1 U3825 ( .A1(n3068), .A2(n3067), .A3(n3066), .A4(n3065), .Z(n3074)
         );
  HDOAI22D1 U3826 ( .A1(n3104), .A2(n1789), .B1(n3103), .B2(n3561), .Z(n3065)
         );
  HDOAI22D1 U3827 ( .A1(n3094), .A2(n3563), .B1(n3093), .B2(n3560), .Z(n3066)
         );
  HDOAI22D1 U3828 ( .A1(n3076), .A2(n1783), .B1(n3075), .B2(n3576), .Z(n3067)
         );
  HDOAI22D1 U3829 ( .A1(n3058), .A2(n2686), .B1(n3057), .B2(n2702), .Z(n3068)
         );
  HDOAI22D1 U3830 ( .A1(n3257), .A2(n2710), .B1(n3179), .B2(n2708), .Z(n3063)
         );
  HDOAI22D1 U3831 ( .A1(n3060), .A2(n2456), .B1(n3111), .B2(n2704), .Z(n3064)
         );
  HDNOR2D1 U3832 ( .A1(n3137), .A2(n2704), .Z(n3090) );
  HDOAI22D1 U3833 ( .A1(n3165), .A2(n3513), .B1(n3553), .B2(n3096), .Z(n3086)
         );
  HDNOR2D1 U3834 ( .A1(n3224), .A2(n2704), .Z(n3087) );
  HDNOR2D1 U3835 ( .A1(n3119), .A2(n2704), .Z(n3082) );
  HDOAI22D1 U3836 ( .A1(n3165), .A2(n3505), .B1(n3394), .B2(n3096), .Z(n3078)
         );
  HDOAI22D1 U3837 ( .A1(n3287), .A2(n2456), .B1(n3203), .B2(n2704), .Z(n3079)
         );
  HDOAI21D1 U3838 ( .A1(n2703), .A2(byp_alu_rs1_data_e[19]), .B(n1769), .Z(
        n3053) );
  HDNOR4D1 U3839 ( .A1(n3050), .A2(n3051), .A3(n3049), .A4(n3048), .Z(n3056)
         );
  HDOAI22D1 U3840 ( .A1(n3094), .A2(n1789), .B1(n3093), .B2(n3561), .Z(n3048)
         );
  HDNAN2D1 U3841 ( .A1(n3045), .A2(ecl_shft_shift4_e[3]), .Z(n3046) );
  HDINVD1 U3842 ( .A(n3240), .Z(n3045) );
  HDAOI22D1 U3843 ( .A1(n3099), .A2(ecl_shft_shift4_e[1]), .B1(n3043), .B2(
        ecl_shft_shift4_e[0]), .Z(n3047) );
  HDAOI22M10D1 U3844 ( .B1(n2680), .B2(n3100), .A1(n2655), .A2(n3336), .Z(
        n2851) );
  HDNAN3D1 U3845 ( .A1(n2909), .A2(n3142), .A3(n2961), .Z(n3099) );
  HDAOI22M10D1 U3846 ( .B1(n2680), .B2(n3159), .A1(n2696), .A2(n3370), .Z(
        n2909) );
  HDOAI22M10D1 U3847 ( .A1(n3237), .A2(n2675), .B1(n3239), .B2(n2655), .Z(
        n2980) );
  HDOAI22D1 U3848 ( .A1(n3340), .A2(n3165), .B1(n3241), .B2(n2456), .Z(n3042)
         );
  HDOAI22D1 U3849 ( .A1(n3076), .A2(n3563), .B1(n3075), .B2(n3560), .Z(n3049)
         );
  HDAOI22D1 U3850 ( .A1(n3092), .A2(ecl_shft_shift4_e[1]), .B1(
        ecl_shft_shift4_e[0]), .B2(n3022), .Z(n3023) );
  HDNAN3D1 U3851 ( .A1(n2833), .A2(n3077), .A3(n2961), .Z(n3022) );
  HDAOI22D1 U3852 ( .A1(n2695), .A2(n3327), .B1(n2682), .B2(n3088), .Z(n2833)
         );
  HDNAN3D1 U3853 ( .A1(n2889), .A2(n3123), .A3(n2961), .Z(n3092) );
  HDNAN2D1 U3854 ( .A1(n3021), .A2(ecl_shft_shift4_e[3]), .Z(n3024) );
  HDINVD1 U3855 ( .A(n3220), .Z(n3021) );
  HDAND3D1 U3856 ( .A1(n3201), .A2(n2961), .A3(n2960), .Z(n3137) );
  HDAOI22M10D1 U3857 ( .B1(n2680), .B2(n3216), .A1(n2299), .A2(n3398), .Z(
        n2960) );
  HDOAI22D1 U3858 ( .A1(n3096), .A2(n3513), .B1(n3553), .B2(n3040), .Z(n3017)
         );
  HDOAI22D1 U3859 ( .A1(n3058), .A2(n1783), .B1(n3057), .B2(n3576), .Z(n3050)
         );
  HDAND3D1 U3860 ( .A1(n2945), .A2(n3182), .A3(n2961), .Z(n3119) );
  HDOAI22D1 U3861 ( .A1(n3320), .A2(n3165), .B1(n3203), .B2(n2456), .Z(n3007)
         );
  HDOAI22D1 U3862 ( .A1(n3038), .A2(n2686), .B1(n3037), .B2(n2702), .Z(n3051)
         );
  HDOAI22D1 U3863 ( .A1(n3179), .A2(n2710), .B1(n3111), .B2(n2708), .Z(n3003)
         );
  HDOAI22D1 U3864 ( .A1(n3060), .A2(n2704), .B1(n2999), .B2(n2456), .Z(n3004)
         );
  HDAND3D1 U3865 ( .A1(n3039), .A2(n2961), .A3(n2803), .Z(n2999) );
  HDAOI22M10D1 U3866 ( .B1(n2681), .B2(n3061), .A1(n2299), .A2(n3311), .Z(
        n2803) );
  HDAOI22M10D1 U3867 ( .B1(n2680), .B2(n3112), .A1(n2655), .A2(n3344), .Z(
        n2868) );
  HDOAI22D1 U3868 ( .A1(n3316), .A2(n3165), .B1(n3184), .B2(n2456), .Z(n2998)
         );
  HDOAI211D1 U3869 ( .A1(ecl_alu_out_sel_shift_e_l), .A2(n3256), .B(n3255), 
        .C(n3254), .Z(alu_byp_rd_data_e[31]) );
  HDAOI22D1 U3870 ( .A1(byp_alu_rs2_data_e[31]), .A2(n2683), .B1(
        alu_adder_out[31]), .B2(n1785), .Z(n3254) );
  HDAOI22D1 U3871 ( .A1(alu_addsub_rs2_data[31]), .A2(n3253), .B1(n3252), .B2(
        byp_alu_rs1_data_e[31]), .Z(n3255) );
  HDOAI211D1 U3872 ( .A1(alu_addsub_rs2_data[31]), .A2(n2703), .B(n1769), .C(
        n3251), .Z(n3252) );
  HDOAI21D1 U3873 ( .A1(n2703), .A2(byp_alu_rs1_data_e[31]), .B(n1769), .Z(
        n3253) );
  HDNOR4D1 U3874 ( .A1(n3250), .A2(n3249), .A3(n3248), .A4(n3247), .Z(n3256)
         );
  HDOAI22D1 U3875 ( .A1(n3292), .A2(n3560), .B1(n3291), .B2(n3563), .Z(n3247)
         );
  HDOAI22D1 U3876 ( .A1(n3246), .A2(n2702), .B1(n3245), .B2(n3533), .Z(n3249)
         );
  HDOAI22D1 U3877 ( .A1(n3257), .A2(n2704), .B1(n3179), .B2(n2456), .Z(n3180)
         );
  HDOAI22D1 U3878 ( .A1(n3345), .A2(n2710), .B1(n3178), .B2(n2708), .Z(n3181)
         );
  HDOAI22D1 U3879 ( .A1(n3294), .A2(n3561), .B1(n3293), .B2(n1789), .Z(n3250)
         );
  HDOAI22D1 U3880 ( .A1(n3374), .A2(n2710), .B1(n3411), .B2(n2707), .Z(n2576)
         );
  HDOAI22D1 U3881 ( .A1(n3443), .A2(n2709), .B1(n3481), .B2(n2710), .Z(n3371)
         );
  HDNOR2D1 U3882 ( .A1(n3408), .A2(n2704), .Z(n3372) );
  HDOAI22D1 U3883 ( .A1(n3421), .A2(n2709), .B1(n3384), .B2(n2710), .Z(n3385)
         );
  HDNAN2M1D1 U3884 ( .A1(n2689), .A2(byp_alu_rs2_data_e[50]), .Z(n2517) );
  HDOAI21D1 U3885 ( .A1(n2703), .A2(byp_alu_rs1_data_e[50]), .B(n1769), .Z(
        n2519) );
  HDNAN3D1 U3886 ( .A1(n1769), .A2(n2520), .A3(n2521), .Z(n2518) );
  HDNAN2D1 U3887 ( .A1(n1772), .A2(n2522), .Z(n2520) );
  HDOAI21D1 U3888 ( .A1(n1994), .A2(n3533), .B(n2526), .Z(n2525) );
  HDOAI22D1 U3889 ( .A1(n3453), .A2(n3560), .B1(n3451), .B2(n3576), .Z(n2527)
         );
  HDOAI22D1 U3890 ( .A1(n3468), .A2(n1789), .B1(n3452), .B2(n3563), .Z(n2523)
         );
  HDOAI22D1 U3891 ( .A1(n3434), .A2(n2705), .B1(n3472), .B2(n2710), .Z(n3365)
         );
  HDNOR2D1 U3892 ( .A1(n3399), .A2(n2704), .Z(n3366) );
  HDOAI22D1 U3893 ( .A1(n3429), .A2(n2709), .B1(n3462), .B2(n2710), .Z(n3352)
         );
  HDNOR2D1 U3894 ( .A1(n3390), .A2(n2704), .Z(n3353) );
  HDOAI22D1 U3895 ( .A1(n2585), .A2(n2707), .B1(n3358), .B2(n2710), .Z(n3359)
         );
  HDNAN2M1D1 U3896 ( .A1(n2689), .A2(byp_alu_rs2_data_e[58]), .Z(n2595) );
  HDOAI21D1 U3897 ( .A1(n2703), .A2(byp_alu_rs1_data_e[58]), .B(n1769), .Z(
        n2597) );
  HDNAN3D1 U3898 ( .A1(n1769), .A2(n2598), .A3(n2599), .Z(n2596) );
  HDNAN2D1 U3899 ( .A1(n1772), .A2(n2600), .Z(n2598) );
  HDOAI21D1 U3900 ( .A1(n3525), .A2(n3563), .B(n2602), .Z(n2601) );
  HDNOR2D1 U3901 ( .A1(n3519), .A2(n3576), .Z(n2605) );
  HDOAI22D1 U3902 ( .A1(n3545), .A2(n3561), .B1(n3526), .B2(n3560), .Z(n2604)
         );
  HDNOR2D1 U3903 ( .A1(n3509), .A2(n2702), .Z(n2603) );
  HDNOR2D1 U3904 ( .A1(n3462), .A2(n2705), .Z(n3391) );
  HDOAI22D1 U3905 ( .A1(n3429), .A2(n2704), .B1(n3390), .B2(n2456), .Z(n3392)
         );
  HDNOR2D1 U3906 ( .A1(n3345), .A2(n2704), .Z(n3312) );
  HDOAI22D1 U3907 ( .A1(n3443), .A2(n2710), .B1(n3408), .B2(n2707), .Z(n3337)
         );
  HDOAI22D1 U3908 ( .A1(n3434), .A2(n2710), .B1(n3399), .B2(n2707), .Z(n3330)
         );
  HDOAI22D1 U3909 ( .A1(n3349), .A2(n2710), .B1(n3384), .B2(n2705), .Z(n3350)
         );
  HDNOR2D1 U3910 ( .A1(n3421), .A2(n2704), .Z(n3351) );
  HDOAI22D1 U3911 ( .A1(n2584), .A2(n2704), .B1(n2510), .B2(n2456), .Z(n3321)
         );
  HDNOR2D1 U3912 ( .A1(n3358), .A2(n2705), .Z(n3322) );
  HDOAI22D1 U3913 ( .A1(n3374), .A2(n2704), .B1(n3411), .B2(n2456), .Z(n3307)
         );
  HDOAI22D1 U3914 ( .A1(n2704), .A2(n3358), .B1(n2584), .B2(n2456), .Z(n3289)
         );
  HDNOR2D1 U3915 ( .A1(n3287), .A2(n2710), .Z(n3290) );
  HDOAI22D1 U3916 ( .A1(n3284), .A2(n2456), .B1(n3319), .B2(n2704), .Z(n3285)
         );
  HDNOR2D1 U3917 ( .A1(n3390), .A2(n2710), .Z(n3286) );
  HDNOR2D1 U3918 ( .A1(n3472), .A2(n2706), .Z(n3400) );
  HDOAI22D1 U3919 ( .A1(n3434), .A2(n2704), .B1(n3399), .B2(n2456), .Z(n3401)
         );
  HDOAI22D1 U3920 ( .A1(n3499), .A2(n2704), .B1(n2106), .B2(n2456), .Z(n3423)
         );
  HDNOR2D1 U3921 ( .A1(n3421), .A2(n2710), .Z(n3424) );
  HDOAI22D1 U3922 ( .A1(n3454), .A2(n2710), .B1(n3493), .B2(n2707), .Z(n3419)
         );
  HDNOR2D1 U3923 ( .A1(n3416), .A2(n2456), .Z(n3420) );
  HDOAI22D1 U3924 ( .A1(n3429), .A2(n2456), .B1(n3462), .B2(n2704), .Z(n3430)
         );
  HDNAN2D1 U3925 ( .A1(n2138), .A2(byp_alu_rs1_data_e[35]), .Z(n3304) );
  HDNOR2D1 U3926 ( .A1(n3481), .A2(n2706), .Z(n3409) );
  HDOAI22D1 U3927 ( .A1(n3443), .A2(n2704), .B1(n3408), .B2(n2456), .Z(n3410)
         );
  HDOAI22D1 U3928 ( .A1(n1877), .A2(n2704), .B1(n2002), .B2(n2456), .Z(n3441)
         );
  HDNOR2D1 U3929 ( .A1(n3478), .A2(n2706), .Z(n3442) );
  HDNAN2D1 U3930 ( .A1(n2699), .A2(byp_alu_rs1_data_e[38]), .Z(n2587) );
  HDOAI22D1 U3931 ( .A1(n3434), .A2(n2456), .B1(n3472), .B2(n2704), .Z(n3435)
         );
  HDOAI22D1 U3932 ( .A1(n3524), .A2(n2704), .B1(n2706), .B2(n2124), .Z(n2512)
         );
  HDOAI22D1 U3933 ( .A1(n3443), .A2(n2456), .B1(n3481), .B2(n2704), .Z(n3444)
         );
  HDOAI211D1 U3934 ( .A1(ecl_alu_out_sel_shift_e_l), .A2(n3281), .B(n3280), 
        .C(n3279), .Z(alu_byp_rd_data_e[32]) );
  HDNAN2D1 U3935 ( .A1(n3275), .A2(n1769), .Z(n3276) );
  HDOAI21D1 U3936 ( .A1(n2703), .A2(byp_alu_rs1_data_e[32]), .B(n1769), .Z(
        n3277) );
  HDNOR4D1 U3937 ( .A1(n3274), .A2(n3273), .A3(n3272), .A4(n3271), .Z(n3281)
         );
  HDOAI22D1 U3938 ( .A1(n3292), .A2(n3576), .B1(n3291), .B2(n1783), .Z(n3271)
         );
  HDINVD1 U3939 ( .A(n3298), .Z(n3223) );
  HDNOR2D1 U3940 ( .A1(n2675), .A2(n3436), .Z(n3014) );
  HDAND2D1 U3941 ( .A1(n1782), .A2(n2786), .Z(n3015) );
  HDOAI22D1 U3942 ( .A1(n3296), .A2(n2704), .B1(n3220), .B2(n2456), .Z(n3221)
         );
  HDOAI22D1 U3943 ( .A1(n3328), .A2(n2708), .B1(n3219), .B2(n2710), .Z(n3222)
         );
  HDNAN2D1 U3944 ( .A1(n1782), .A2(n3216), .Z(n3217) );
  HDINVD1 U3945 ( .A(n3398), .Z(n3218) );
  HDOAI22D1 U3946 ( .A1(n3294), .A2(n3560), .B1(n3293), .B2(n3563), .Z(n3272)
         );
  HDINVD1 U3947 ( .A(n3567), .Z(n3000) );
  HDNOR2D1 U3948 ( .A1(n3241), .A2(n2710), .Z(n3244) );
  HDNAN2D1 U3949 ( .A1(n2203), .A2(byp_alu_rs1_data_e[19]), .Z(n3039) );
  HDOA21D1 U3950 ( .A1(n3431), .A2(n2675), .B(n3005), .Z(n3203) );
  HDNAN2D1 U3951 ( .A1(n2662), .A2(byp_alu_rs1_data_e[21]), .Z(n3077) );
  HDINVD1 U3952 ( .A(n3354), .Z(n3199) );
  HDNAN2D1 U3953 ( .A1(n1782), .A2(n3196), .Z(n3197) );
  HDOAI22D1 U3954 ( .A1(n3349), .A2(n2704), .B1(n3384), .B2(n2456), .Z(n3267)
         );
  HDNAN2D1 U3955 ( .A1(n2699), .A2(byp_alu_rs1_data_e[28]), .Z(n3182) );
  HDNOR2D1 U3956 ( .A1(n3264), .A2(n2710), .Z(n3268) );
  HDNAN2D1 U3957 ( .A1(n2701), .A2(byp_alu_rs1_data_e[24]), .Z(n3107) );
  HDOAI22D1 U3958 ( .A1(n3378), .A2(n2710), .B1(n3345), .B2(n2705), .Z(n3262)
         );
  HDOAI211D1 U3959 ( .A1(n3114), .A2(n2109), .B(n3260), .C(n3113), .Z(n3314)
         );
  HDINVD1 U3960 ( .A(n3344), .Z(n3114) );
  HDAOI22D1 U3961 ( .A1(n2609), .A2(alu_addsub_rs2_data[62]), .B1(n2610), .B2(
        byp_alu_rs1_data_e[62]), .Z(n2608) );
  HDOAI211D1 U3962 ( .A1(n2703), .A2(alu_addsub_rs2_data[62]), .B(n1769), .C(
        n2611), .Z(n2610) );
  HDNAN2D1 U3963 ( .A1(n1767), .A2(alu_addsub_rs2_data[62]), .Z(n2611) );
  HDOAI21D1 U3964 ( .A1(n2703), .A2(byp_alu_rs1_data_e[62]), .B(n1769), .Z(
        n2609) );
  HDNAN4M2D1 U3965 ( .A1(n2613), .A2(n3577), .A3(n2614), .A4(n2615), .Z(n2612)
         );
  HDOAI22D1 U3966 ( .A1(n3540), .A2(n2705), .B1(n3539), .B2(n2710), .Z(n3541)
         );
  HDAOI21D1 U3967 ( .A1(n3538), .A2(n3537), .B(n2456), .Z(n3542) );
  HDOAI211D1 U3968 ( .A1(n2002), .A2(n2710), .B(n3558), .C(n3557), .Z(n3571)
         );
  HDAOI22D1 U3969 ( .A1(n3555), .A2(ecl_shft_shift4_e[0]), .B1(n3554), .B2(
        ecl_shft_shift4_e[1]), .Z(n3558) );
  HDOAI211D1 U3970 ( .A1(n3553), .A2(n2008), .B(n3552), .C(n3551), .Z(n3555)
         );
  HDAOI22D1 U3971 ( .A1(n3550), .A2(byp_alu_rs1_data_e[30]), .B1(n2691), .B2(
        byp_alu_rs1_data_e[46]), .Z(n3551) );
  HDAOI211D1 U3972 ( .A1(n2651), .A2(n1924), .B(n2650), .C(n2652), .Z(n2643)
         );
  HDINVD1 U3973 ( .A(alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_28_), .Z(
        n2645) );
  HDAOI21M10D1 U3974 ( .A1(n3526), .A2(n2503), .B(n2647), .Z(n2646) );
  HDOAI222D1 U3975 ( .A1(n3564), .A2(n3560), .B1(n3574), .B2(n3561), .C1(n3545), .C2(n3576), .Z(n2647) );
  HDAOI21D1 U3976 ( .A1(n3510), .A2(ecl_shft_shift4_e[0]), .B(n3527), .Z(n3545) );
  HDAOI21D1 U3977 ( .A1(n3520), .A2(ecl_shft_shift4_e[0]), .B(n3527), .Z(n3564) );
  HDOR2D1 U3978 ( .A1(n3544), .A2(n3563), .Z(n2649) );
  HDAOI22M10D1 U3979 ( .B1(n2502), .B2(ecl_shft_shift4_e[0]), .A1(n2704), .A2(
        n3570), .Z(n3522) );
  HDOAI211D1 U3980 ( .A1(n3521), .A2(n2008), .B(n2546), .C(n2545), .Z(n2502)
         );
  HDAOI22D1 U3981 ( .A1(n3550), .A2(byp_alu_rs1_data_e[27]), .B1(n2691), .B2(
        byp_alu_rs1_data_e[43]), .Z(n2546) );
  HDOA222D1 U3982 ( .A1(n2106), .A2(n2710), .B1(n2547), .B2(n2456), .C1(n3531), 
        .C2(n2705), .Z(n2550) );
  HDAOI211D1 U3983 ( .A1(n2691), .A2(byp_alu_rs1_data_e[44]), .B(n2548), .C(
        n2549), .Z(n2547) );
  HDOAI22D1 U3984 ( .A1(n1877), .A2(n2710), .B1(n2002), .B2(n2708), .Z(n3517)
         );
  HDOAI211D1 U3985 ( .A1(n3513), .A2(n2008), .B(n3512), .C(n3511), .Z(n3554)
         );
  HDAOI22D1 U3986 ( .A1(n3550), .A2(byp_alu_rs1_data_e[26]), .B1(n2691), .B2(
        byp_alu_rs1_data_e[42]), .Z(n3511) );
  HDNAN2D1 U3987 ( .A1(n2698), .A2(byp_alu_rs1_data_e[58]), .Z(n3512) );
  HDOAI22D1 U3988 ( .A1(n3454), .A2(n2709), .B1(n3493), .B2(n2704), .Z(n3455)
         );
  HDOAI22D1 U3989 ( .A1(n3540), .A2(n2456), .B1(n3539), .B2(n2704), .Z(n2619)
         );
  HDNOR2D1 U3990 ( .A1(n3462), .A2(n2456), .Z(n3463) );
  HDNAN2D1 U3991 ( .A1(n2701), .A2(byp_alu_rs1_data_e[42]), .Z(n3363) );
  HDNAN2D1 U3992 ( .A1(n3550), .A2(byp_alu_rs1_data_e[22]), .Z(n3476) );
  HDNAN2D1 U3993 ( .A1(n2138), .A2(byp_alu_rs1_data_e[44]), .Z(n3382) );
  HDAOI22D1 U3994 ( .A1(n3536), .A2(n3458), .B1(n2699), .B2(
        byp_alu_rs1_data_e[52]), .Z(n3459) );
  HDOAI211D1 U3995 ( .A1(n3498), .A2(n2008), .B(n3497), .C(n3496), .Z(n3532)
         );
  HDAOI22D1 U3996 ( .A1(n3550), .A2(byp_alu_rs1_data_e[24]), .B1(n2691), .B2(
        byp_alu_rs1_data_e[40]), .Z(n3496) );
  HDOAI22D1 U3997 ( .A1(n3524), .A2(n2705), .B1(n2124), .B2(n2710), .Z(n3489)
         );
  HDNAN2D1 U3998 ( .A1(n2743), .A2(byp_alu_rs1_data_e[31]), .Z(n3567) );
  HDNOR2D1 U3999 ( .A1(n3481), .A2(n2456), .Z(n3482) );
  HDNOR2D1 U4000 ( .A1(n3540), .A2(n2704), .Z(n3507) );
  HDAOI22D1 U4001 ( .A1(n3550), .A2(byp_alu_rs1_data_e[21]), .B1(n2105), .B2(
        byp_alu_rs1_data_e[37]), .Z(n3466) );
  HDOAI211D1 U4002 ( .A1(n3505), .A2(n2008), .B(n3504), .C(n3503), .Z(n3543)
         );
  HDAOI22D1 U4003 ( .A1(n3550), .A2(byp_alu_rs1_data_e[25]), .B1(n2691), .B2(
        byp_alu_rs1_data_e[41]), .Z(n3503) );
  HDAOI21D1 U4004 ( .A1(n3502), .A2(ecl_shft_shift4_e[0]), .B(n3527), .Z(n3526) );
  HDEXOR2D1 U4005 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[54]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_22_) );
  HDEXOR2D1 U4006 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[53]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_21_) );
  HDEXOR2D1 U4007 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[49]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_17_) );
  HDEXOR2D1 U4008 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[47]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_15_) );
  HDEXOR2D1 U4009 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[46]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_14_) );
  HDEXOR2D1 U4010 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[45]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_13_) );
  HDEXOR2D1 U4011 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[39]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_7_) );
  HDEXOR2D1 U4012 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[37]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_5_) );
  HDEXOR2D1 U4013 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[35]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_3_) );
  HDEXOR2D1 U4014 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[34]), .Z(
        alu_addsub_rs2_data[34]) );
  HDEXOR2D1 U4015 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[30]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I2_30_) );
  HDEXOR2D1 U4016 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[29]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I2_29_) );
  HDEXOR2D1 U4017 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[22]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I2_22_) );
  HDEXOR2D1 U4018 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[20]), .Z(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I2_20_) );
  HDEXOR2D1 U4019 ( .A1(ifu_exu_invert_d), .A2(byp_alu_rs2_data_e[14]), .Z(
        alu_addsub_rs2_data[14]) );
  HDNAN2D1 U4020 ( .A1(n1767), .A2(
        alu_addsub_adder_add_24_2_DP_OP_282_4997_7_I5_28_), .Z(n2644) );
  HDMUXB2DL U4021 ( .A0(n1772), .A1(n1767), .SL(n2146), .Z(n2988) );
  HDMUXB2DL U4022 ( .A0(n1772), .A1(n1767), .SL(alu_addsub_rs2_data[0]), .Z(
        n2758) );
  HDMUXB2DL U4023 ( .A0(n1772), .A1(n1767), .SL(n2007), .Z(n3129) );
  HDMUXB2DL U4024 ( .A0(n1772), .A1(n1767), .SL(alu_addsub_rs2_data[13]), .Z(
        n2951) );
  HDMUXB2DL U4025 ( .A0(n1772), .A1(n1767), .SL(n2176), .Z(n2768) );
  HDMUXB2DL U4026 ( .A0(n1772), .A1(n1767), .SL(n2169), .Z(n2935) );
  HDMUXB2DL U4027 ( .A0(n1772), .A1(n1767), .SL(n2175), .Z(n2971) );
  HDMUXB2DL U4028 ( .A0(n1772), .A1(n1767), .SL(n2173), .Z(n2917) );
  HDMUXB2DL U4029 ( .A0(n1772), .A1(n1767), .SL(n2117), .Z(n3150) );
  HDMUXB2DL U4030 ( .A0(n1772), .A1(n1767), .SL(n2160), .Z(n2826) );
  HDMUXB2DL U4031 ( .A0(n1772), .A1(n1767), .SL(n1880), .Z(n2842) );
  HDMUXB2DL U4032 ( .A0(n1772), .A1(n1767), .SL(n2189), .Z(n2875) );
  HDMUXB2DL U4033 ( .A0(n1772), .A1(n1767), .SL(n2197), .Z(n2858) );
  HDMUXB2DL U4034 ( .A0(n1772), .A1(n1767), .SL(n2171), .Z(n3069) );
  HDMUXB2DL U4035 ( .A0(n1772), .A1(n1767), .SL(n1867), .Z(n3169) );
  HDMUXB2DL U4036 ( .A0(n1772), .A1(n1767), .SL(n1979), .Z(n3231) );
  HDMUXB2DL U4037 ( .A0(n1772), .A1(n1767), .SL(n1976), .Z(n3190) );
  HDMUXB2DL U4038 ( .A0(n1772), .A1(n1767), .SL(n1969), .Z(n3210) );
  HDMUXB2DL U4039 ( .A0(n1772), .A1(n1767), .SL(n2148), .Z(n3031) );
  HDMUXB2DL U4040 ( .A0(n1772), .A1(n1767), .SL(n2137), .Z(n3275) );
endmodule

